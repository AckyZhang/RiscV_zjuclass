`timescale 1ns/100ps
//correct read result:
// 000004dd 000006c4 000006de 000003bb 000006db 000006d7 0000027c 00000278 00000628 00000646 00000590 0000039d 00000472 00000780 000001a3 00000031 0000000e 00000266 00000578 000003e1 000003c4 00000377 00000288 000001e2 00000224 000001da 00000765 000006c4 0000036b 00000753 00000058 00000526 000004be 000003a5 0000045a 000003bb 0000068a 00000547 000002af 00000533 000000af 00000290 00000688 00000654 00000771 0000011a 00000012 000007c2 0000007c 000000b5 0000011f 000003d8 0000061a 000003d0 000000c2 000002af 0000055f 00000763 000001aa 000003d7 000000be 00000767 000007e9 00000741 000000a9 0000069a 00000406 00000083 0000012f 00000316 000004a9 000006b1 000002bb 000001fb 0000053f 0000033b 00000002 0000011d 0000061a 0000005d 000003fc 000004a6 000001cb 00000273 000003b1 00000084 000000e2 00000089 00000519 0000044e 000004cf 000001f5 000004c0 00000312 00000049 000002ba 0000074e 00000390 0000065e 000000c8 0000008e 0000015b 000006a7 000000da 0000029d 00000281 000004eb 00000704 000007aa 0000022e 000004c5 00000241 00000071 000003b4 00000534 0000042d 000000a0 00000488 000000f2 00000170 00000441 0000004d 00000514 00000781 000007f0 0000074b 000004eb 0000024f 000002c9 000002c1 0000028e 00000549 000001af 000001d5 000003ad 00000635 0000018c 000006e5 00000432 00000530 0000019e 00000588 000003c9 0000043d 0000061e 0000023a 000000aa 00000203 0000056f 000004b5 000002b2 000002e3 000007d9 000001c6 00000290 000002e7 000001f9 000001dd 00000041 000001e1 00000402 000002bd 000004b9 00000595 00000740 000002be 00000699 0000073d 0000020d 0000024b 0000059e 0000035f 00000241 00000288 00000479 000002b4 000000a9 00000555 000002f7 0000003b 0000067b 000002b4 00000327 0000012a 000001a6 000005cf 000000da 0000025d 0000018d 000003c5 0000078b 00000215 0000033e 0000068a 0000076c 00000712 00000589 00000778 000003fa 00000546 000002d9 000005e8 0000059d 00000235 000003cb 000002ba 00000670 00000150 0000077a 00000530 0000070a 00000143 000006e7 00000116 0000031d 000007e1 000005dd 00000031 000003bf 0000051a 000006e8 00000244 000000a5 000005e4 00000597 000004c0 000006cb 000007ca 0000014f 00000555 000003d0 00000374 0000046a 00000344 00000111 00000210 000007a3 0000001d 00000587 000002a5 0000042a 000000d6 000003d3 0000072e 000004d6 0000001e 00000677 0000007b 0000044a 000007d1 00000224 00000210 0000011f 000005ed 00000243 00000223 00000382 00000453 00000050 000001db 00000227 000001c2 000005df 000002ac 00000595 00000057 0000029a 000003f7 00000068 000003aa 000006cf 00000029 000004c3 0000057d 00000791 0000076c 000005fe 00000273 00000153 000004f4 00000691 000003fc 0000028b 0000008f 000006d9 00000024 0000034c 00000628 000003d5 0000065d 000006fa 000006a9 00000170 00000094 00000431 000007ca 00000438 0000063d 0000071b 00000184 000005a5 00000096 0000026f 00000591 0000004e 00000034 0000020c 000001dc 000000bb 0000079f 0000064e 00000693 00000484 00000618 00000776 00000403 000005f6 00000302 000005b1 000004a9 000007e9 000000b8 000006a6 00000726 000002a8 00000438 000001d1 000006fa 0000035b 000000de 000000e4 00000617 000003b1 00000166 00000498 000007e0 0000020c 00000542 00000106 00000559 000003cb 00000366 0000017b 00000750 00000735 000003f2 0000017b 000007e9 000001d3 0000054e 00000098 00000081 00000103 00000547 000006b7 000001b7 00000542 00000729 0000055e 000002ea 00000527 000007d2 000004ed 00000225 000002e9 00000266 00000339 00000277 00000163 0000071d 000007b9 000006a6 00000705 00000553 000000a3 0000062c 00000279 000006f4 00000548 00000313 000005c2 000001b0 000002e7 000000b9 0000033c 000003c7 0000056d 000004bb 00000665 00000115 00000391 0000027b 00000468 000004fc 00000005 000003e1 00000526 000000f1 000002cc 000007e9 0000011f 000004a0 0000072b 0000026f 0000008c 000004ec 00000149 00000248 000001da 000006f8 000002ae 000003a3 0000025f 00000761 00000000 000005e0 000002f5 000001d8 00000225 0000040c 000007a7 00000521 00000617 00000664 000002d3 0000040a 00000398 00000463 00000240 0000018a 000007ad 0000043d 00000487 0000062e 00000003 00000431 000000c3 00000153 000003e1 000000c1 000002a7 0000010e 000001f5 00000396 00000589 00000605 00000307 00000123 00000581 00000527 0000050b 0000038e 00000092 000002ac 000002e1 0000053b 0000062c 000000b6 0000054e 0000027a 000000d7 00000669 0000052e 000002eb 000004db 00000526 00000704 00000508 000004d5 00000690 00000387 00000556 00000398 0000049b 00000640 000004a2 0000003d 000005fd 00000525 000003aa 00000348 000001c8 000000d1 00000479 000002f5 0000044f 000003a3 0000039c 00000175 000001e7 000003e1 000001fc 000003b0 000005ad 00000362 0000061e 00000690 000000da 0000079e 000007fd 000000ea 000006ea 0000028f 00000379 0000073a 00000666 00000500 00000628 00000035 000007d6 000007e2 00000694

module cache_tb();

`define DATA_COUNT (512)
`define RDWR_COUNT (6*`DATA_COUNT)

reg wr_cycle           [`RDWR_COUNT];
reg rd_cycle           [`RDWR_COUNT];
reg [31:0] addr_rom    [`RDWR_COUNT];
reg [31:0] wr_data_rom [`RDWR_COUNT];
reg [31:0] validation_data [`DATA_COUNT];

initial begin
    // 512 sequence write cycles
    rd_cycle[    0] = 1'b0;  wr_cycle[    0] = 1'b1;  addr_rom[    0]='h00000000;  wr_data_rom[    0]='h00000114;
    rd_cycle[    1] = 1'b0;  wr_cycle[    1] = 1'b1;  addr_rom[    1]='h00000004;  wr_data_rom[    1]='h00000728;
    rd_cycle[    2] = 1'b0;  wr_cycle[    2] = 1'b1;  addr_rom[    2]='h00000008;  wr_data_rom[    2]='h000006de;
    rd_cycle[    3] = 1'b0;  wr_cycle[    3] = 1'b1;  addr_rom[    3]='h0000000c;  wr_data_rom[    3]='h000006cd;
    rd_cycle[    4] = 1'b0;  wr_cycle[    4] = 1'b1;  addr_rom[    4]='h00000010;  wr_data_rom[    4]='h000006cf;
    rd_cycle[    5] = 1'b0;  wr_cycle[    5] = 1'b1;  addr_rom[    5]='h00000014;  wr_data_rom[    5]='h000002d4;
    rd_cycle[    6] = 1'b0;  wr_cycle[    6] = 1'b1;  addr_rom[    6]='h00000018;  wr_data_rom[    6]='h00000452;
    rd_cycle[    7] = 1'b0;  wr_cycle[    7] = 1'b1;  addr_rom[    7]='h0000001c;  wr_data_rom[    7]='h000002d7;
    rd_cycle[    8] = 1'b0;  wr_cycle[    8] = 1'b1;  addr_rom[    8]='h00000020;  wr_data_rom[    8]='h00000130;
    rd_cycle[    9] = 1'b0;  wr_cycle[    9] = 1'b1;  addr_rom[    9]='h00000024;  wr_data_rom[    9]='h00000745;
    rd_cycle[   10] = 1'b0;  wr_cycle[   10] = 1'b1;  addr_rom[   10]='h00000028;  wr_data_rom[   10]='h00000253;
    rd_cycle[   11] = 1'b0;  wr_cycle[   11] = 1'b1;  addr_rom[   11]='h0000002c;  wr_data_rom[   11]='h00000494;
    rd_cycle[   12] = 1'b0;  wr_cycle[   12] = 1'b1;  addr_rom[   12]='h00000030;  wr_data_rom[   12]='h00000472;
    rd_cycle[   13] = 1'b0;  wr_cycle[   13] = 1'b1;  addr_rom[   13]='h00000034;  wr_data_rom[   13]='h0000006e;
    rd_cycle[   14] = 1'b0;  wr_cycle[   14] = 1'b1;  addr_rom[   14]='h00000038;  wr_data_rom[   14]='h00000096;
    rd_cycle[   15] = 1'b0;  wr_cycle[   15] = 1'b1;  addr_rom[   15]='h0000003c;  wr_data_rom[   15]='h000005ed;
    rd_cycle[   16] = 1'b0;  wr_cycle[   16] = 1'b1;  addr_rom[   16]='h00000040;  wr_data_rom[   16]='h0000000e;
    rd_cycle[   17] = 1'b0;  wr_cycle[   17] = 1'b1;  addr_rom[   17]='h00000044;  wr_data_rom[   17]='h000005a3;
    rd_cycle[   18] = 1'b0;  wr_cycle[   18] = 1'b1;  addr_rom[   18]='h00000048;  wr_data_rom[   18]='h00000105;
    rd_cycle[   19] = 1'b0;  wr_cycle[   19] = 1'b1;  addr_rom[   19]='h0000004c;  wr_data_rom[   19]='h00000465;
    rd_cycle[   20] = 1'b0;  wr_cycle[   20] = 1'b1;  addr_rom[   20]='h00000050;  wr_data_rom[   20]='h00000061;
    rd_cycle[   21] = 1'b0;  wr_cycle[   21] = 1'b1;  addr_rom[   21]='h00000054;  wr_data_rom[   21]='h000003b5;
    rd_cycle[   22] = 1'b0;  wr_cycle[   22] = 1'b1;  addr_rom[   22]='h00000058;  wr_data_rom[   22]='h000005d2;
    rd_cycle[   23] = 1'b0;  wr_cycle[   23] = 1'b1;  addr_rom[   23]='h0000005c;  wr_data_rom[   23]='h00000553;
    rd_cycle[   24] = 1'b0;  wr_cycle[   24] = 1'b1;  addr_rom[   24]='h00000060;  wr_data_rom[   24]='h00000021;
    rd_cycle[   25] = 1'b0;  wr_cycle[   25] = 1'b1;  addr_rom[   25]='h00000064;  wr_data_rom[   25]='h000001da;
    rd_cycle[   26] = 1'b0;  wr_cycle[   26] = 1'b1;  addr_rom[   26]='h00000068;  wr_data_rom[   26]='h000005b7;
    rd_cycle[   27] = 1'b0;  wr_cycle[   27] = 1'b1;  addr_rom[   27]='h0000006c;  wr_data_rom[   27]='h0000051b;
    rd_cycle[   28] = 1'b0;  wr_cycle[   28] = 1'b1;  addr_rom[   28]='h00000070;  wr_data_rom[   28]='h000002b0;
    rd_cycle[   29] = 1'b0;  wr_cycle[   29] = 1'b1;  addr_rom[   29]='h00000074;  wr_data_rom[   29]='h000007b1;
    rd_cycle[   30] = 1'b0;  wr_cycle[   30] = 1'b1;  addr_rom[   30]='h00000078;  wr_data_rom[   30]='h00000037;
    rd_cycle[   31] = 1'b0;  wr_cycle[   31] = 1'b1;  addr_rom[   31]='h0000007c;  wr_data_rom[   31]='h000006d5;
    rd_cycle[   32] = 1'b0;  wr_cycle[   32] = 1'b1;  addr_rom[   32]='h00000080;  wr_data_rom[   32]='h000002f3;
    rd_cycle[   33] = 1'b0;  wr_cycle[   33] = 1'b1;  addr_rom[   33]='h00000084;  wr_data_rom[   33]='h0000021b;
    rd_cycle[   34] = 1'b0;  wr_cycle[   34] = 1'b1;  addr_rom[   34]='h00000088;  wr_data_rom[   34]='h00000584;
    rd_cycle[   35] = 1'b0;  wr_cycle[   35] = 1'b1;  addr_rom[   35]='h0000008c;  wr_data_rom[   35]='h000000ed;
    rd_cycle[   36] = 1'b0;  wr_cycle[   36] = 1'b1;  addr_rom[   36]='h00000090;  wr_data_rom[   36]='h000005d9;
    rd_cycle[   37] = 1'b0;  wr_cycle[   37] = 1'b1;  addr_rom[   37]='h00000094;  wr_data_rom[   37]='h000006a8;
    rd_cycle[   38] = 1'b0;  wr_cycle[   38] = 1'b1;  addr_rom[   38]='h00000098;  wr_data_rom[   38]='h00000360;
    rd_cycle[   39] = 1'b0;  wr_cycle[   39] = 1'b1;  addr_rom[   39]='h0000009c;  wr_data_rom[   39]='h000005b4;
    rd_cycle[   40] = 1'b0;  wr_cycle[   40] = 1'b1;  addr_rom[   40]='h000000a0;  wr_data_rom[   40]='h000000af;
    rd_cycle[   41] = 1'b0;  wr_cycle[   41] = 1'b1;  addr_rom[   41]='h000000a4;  wr_data_rom[   41]='h00000327;
    rd_cycle[   42] = 1'b0;  wr_cycle[   42] = 1'b1;  addr_rom[   42]='h000000a8;  wr_data_rom[   42]='h00000688;
    rd_cycle[   43] = 1'b0;  wr_cycle[   43] = 1'b1;  addr_rom[   43]='h000000ac;  wr_data_rom[   43]='h00000724;
    rd_cycle[   44] = 1'b0;  wr_cycle[   44] = 1'b1;  addr_rom[   44]='h000000b0;  wr_data_rom[   44]='h00000771;
    rd_cycle[   45] = 1'b0;  wr_cycle[   45] = 1'b1;  addr_rom[   45]='h000000b4;  wr_data_rom[   45]='h000001b5;
    rd_cycle[   46] = 1'b0;  wr_cycle[   46] = 1'b1;  addr_rom[   46]='h000000b8;  wr_data_rom[   46]='h00000350;
    rd_cycle[   47] = 1'b0;  wr_cycle[   47] = 1'b1;  addr_rom[   47]='h000000bc;  wr_data_rom[   47]='h0000031c;
    rd_cycle[   48] = 1'b0;  wr_cycle[   48] = 1'b1;  addr_rom[   48]='h000000c0;  wr_data_rom[   48]='h0000007c;
    rd_cycle[   49] = 1'b0;  wr_cycle[   49] = 1'b1;  addr_rom[   49]='h000000c4;  wr_data_rom[   49]='h0000030f;
    rd_cycle[   50] = 1'b0;  wr_cycle[   50] = 1'b1;  addr_rom[   50]='h000000c8;  wr_data_rom[   50]='h000004c9;
    rd_cycle[   51] = 1'b0;  wr_cycle[   51] = 1'b1;  addr_rom[   51]='h000000cc;  wr_data_rom[   51]='h000003d8;
    rd_cycle[   52] = 1'b0;  wr_cycle[   52] = 1'b1;  addr_rom[   52]='h000000d0;  wr_data_rom[   52]='h00000372;
    rd_cycle[   53] = 1'b0;  wr_cycle[   53] = 1'b1;  addr_rom[   53]='h000000d4;  wr_data_rom[   53]='h00000320;
    rd_cycle[   54] = 1'b0;  wr_cycle[   54] = 1'b1;  addr_rom[   54]='h000000d8;  wr_data_rom[   54]='h000000c2;
    rd_cycle[   55] = 1'b0;  wr_cycle[   55] = 1'b1;  addr_rom[   55]='h000000dc;  wr_data_rom[   55]='h00000368;
    rd_cycle[   56] = 1'b0;  wr_cycle[   56] = 1'b1;  addr_rom[   56]='h000000e0;  wr_data_rom[   56]='h000007d9;
    rd_cycle[   57] = 1'b0;  wr_cycle[   57] = 1'b1;  addr_rom[   57]='h000000e4;  wr_data_rom[   57]='h000002a1;
    rd_cycle[   58] = 1'b0;  wr_cycle[   58] = 1'b1;  addr_rom[   58]='h000000e8;  wr_data_rom[   58]='h00000770;
    rd_cycle[   59] = 1'b0;  wr_cycle[   59] = 1'b1;  addr_rom[   59]='h000000ec;  wr_data_rom[   59]='h00000641;
    rd_cycle[   60] = 1'b0;  wr_cycle[   60] = 1'b1;  addr_rom[   60]='h000000f0;  wr_data_rom[   60]='h000004f0;
    rd_cycle[   61] = 1'b0;  wr_cycle[   61] = 1'b1;  addr_rom[   61]='h000000f4;  wr_data_rom[   61]='h0000037f;
    rd_cycle[   62] = 1'b0;  wr_cycle[   62] = 1'b1;  addr_rom[   62]='h000000f8;  wr_data_rom[   62]='h00000157;
    rd_cycle[   63] = 1'b0;  wr_cycle[   63] = 1'b1;  addr_rom[   63]='h000000fc;  wr_data_rom[   63]='h00000033;
    rd_cycle[   64] = 1'b0;  wr_cycle[   64] = 1'b1;  addr_rom[   64]='h00000100;  wr_data_rom[   64]='h00000316;
    rd_cycle[   65] = 1'b0;  wr_cycle[   65] = 1'b1;  addr_rom[   65]='h00000104;  wr_data_rom[   65]='h000004db;
    rd_cycle[   66] = 1'b0;  wr_cycle[   66] = 1'b1;  addr_rom[   66]='h00000108;  wr_data_rom[   66]='h00000190;
    rd_cycle[   67] = 1'b0;  wr_cycle[   67] = 1'b1;  addr_rom[   67]='h0000010c;  wr_data_rom[   67]='h00000568;
    rd_cycle[   68] = 1'b0;  wr_cycle[   68] = 1'b1;  addr_rom[   68]='h00000110;  wr_data_rom[   68]='h0000056b;
    rd_cycle[   69] = 1'b0;  wr_cycle[   69] = 1'b1;  addr_rom[   69]='h00000114;  wr_data_rom[   69]='h00000203;
    rd_cycle[   70] = 1'b0;  wr_cycle[   70] = 1'b1;  addr_rom[   70]='h00000118;  wr_data_rom[   70]='h00000467;
    rd_cycle[   71] = 1'b0;  wr_cycle[   71] = 1'b1;  addr_rom[   71]='h0000011c;  wr_data_rom[   71]='h000002f9;
    rd_cycle[   72] = 1'b0;  wr_cycle[   72] = 1'b1;  addr_rom[   72]='h00000120;  wr_data_rom[   72]='h00000614;
    rd_cycle[   73] = 1'b0;  wr_cycle[   73] = 1'b1;  addr_rom[   73]='h00000124;  wr_data_rom[   73]='h000005e7;
    rd_cycle[   74] = 1'b0;  wr_cycle[   74] = 1'b1;  addr_rom[   74]='h00000128;  wr_data_rom[   74]='h0000044b;
    rd_cycle[   75] = 1'b0;  wr_cycle[   75] = 1'b1;  addr_rom[   75]='h0000012c;  wr_data_rom[   75]='h000003a7;
    rd_cycle[   76] = 1'b0;  wr_cycle[   76] = 1'b1;  addr_rom[   76]='h00000130;  wr_data_rom[   76]='h00000539;
    rd_cycle[   77] = 1'b0;  wr_cycle[   77] = 1'b1;  addr_rom[   77]='h00000134;  wr_data_rom[   77]='h00000512;
    rd_cycle[   78] = 1'b0;  wr_cycle[   78] = 1'b1;  addr_rom[   78]='h00000138;  wr_data_rom[   78]='h0000009f;
    rd_cycle[   79] = 1'b0;  wr_cycle[   79] = 1'b1;  addr_rom[   79]='h0000013c;  wr_data_rom[   79]='h000007e9;
    rd_cycle[   80] = 1'b0;  wr_cycle[   80] = 1'b1;  addr_rom[   80]='h00000140;  wr_data_rom[   80]='h000003fc;
    rd_cycle[   81] = 1'b0;  wr_cycle[   81] = 1'b1;  addr_rom[   81]='h00000144;  wr_data_rom[   81]='h0000061a;
    rd_cycle[   82] = 1'b0;  wr_cycle[   82] = 1'b1;  addr_rom[   82]='h00000148;  wr_data_rom[   82]='h00000283;
    rd_cycle[   83] = 1'b0;  wr_cycle[   83] = 1'b1;  addr_rom[   83]='h0000014c;  wr_data_rom[   83]='h000002e8;
    rd_cycle[   84] = 1'b0;  wr_cycle[   84] = 1'b1;  addr_rom[   84]='h00000150;  wr_data_rom[   84]='h000003dd;
    rd_cycle[   85] = 1'b0;  wr_cycle[   85] = 1'b1;  addr_rom[   85]='h00000154;  wr_data_rom[   85]='h0000012a;
    rd_cycle[   86] = 1'b0;  wr_cycle[   86] = 1'b1;  addr_rom[   86]='h00000158;  wr_data_rom[   86]='h000000cc;
    rd_cycle[   87] = 1'b0;  wr_cycle[   87] = 1'b1;  addr_rom[   87]='h0000015c;  wr_data_rom[   87]='h0000040f;
    rd_cycle[   88] = 1'b0;  wr_cycle[   88] = 1'b1;  addr_rom[   88]='h00000160;  wr_data_rom[   88]='h0000051d;
    rd_cycle[   89] = 1'b0;  wr_cycle[   89] = 1'b1;  addr_rom[   89]='h00000164;  wr_data_rom[   89]='h000000c8;
    rd_cycle[   90] = 1'b0;  wr_cycle[   90] = 1'b1;  addr_rom[   90]='h00000168;  wr_data_rom[   90]='h000004ff;
    rd_cycle[   91] = 1'b0;  wr_cycle[   91] = 1'b1;  addr_rom[   91]='h0000016c;  wr_data_rom[   91]='h000001f5;
    rd_cycle[   92] = 1'b0;  wr_cycle[   92] = 1'b1;  addr_rom[   92]='h00000170;  wr_data_rom[   92]='h0000067a;
    rd_cycle[   93] = 1'b0;  wr_cycle[   93] = 1'b1;  addr_rom[   93]='h00000174;  wr_data_rom[   93]='h00000101;
    rd_cycle[   94] = 1'b0;  wr_cycle[   94] = 1'b1;  addr_rom[   94]='h00000178;  wr_data_rom[   94]='h00000049;
    rd_cycle[   95] = 1'b0;  wr_cycle[   95] = 1'b1;  addr_rom[   95]='h0000017c;  wr_data_rom[   95]='h000002ba;
    rd_cycle[   96] = 1'b0;  wr_cycle[   96] = 1'b1;  addr_rom[   96]='h00000180;  wr_data_rom[   96]='h000006ca;
    rd_cycle[   97] = 1'b0;  wr_cycle[   97] = 1'b1;  addr_rom[   97]='h00000184;  wr_data_rom[   97]='h0000061a;
    rd_cycle[   98] = 1'b0;  wr_cycle[   98] = 1'b1;  addr_rom[   98]='h00000188;  wr_data_rom[   98]='h00000345;
    rd_cycle[   99] = 1'b0;  wr_cycle[   99] = 1'b1;  addr_rom[   99]='h0000018c;  wr_data_rom[   99]='h000000c8;
    rd_cycle[  100] = 1'b0;  wr_cycle[  100] = 1'b1;  addr_rom[  100]='h00000190;  wr_data_rom[  100]='h00000356;
    rd_cycle[  101] = 1'b0;  wr_cycle[  101] = 1'b1;  addr_rom[  101]='h00000194;  wr_data_rom[  101]='h00000228;
    rd_cycle[  102] = 1'b0;  wr_cycle[  102] = 1'b1;  addr_rom[  102]='h00000198;  wr_data_rom[  102]='h000006a7;
    rd_cycle[  103] = 1'b0;  wr_cycle[  103] = 1'b1;  addr_rom[  103]='h0000019c;  wr_data_rom[  103]='h000003b8;
    rd_cycle[  104] = 1'b0;  wr_cycle[  104] = 1'b1;  addr_rom[  104]='h000001a0;  wr_data_rom[  104]='h000000d0;
    rd_cycle[  105] = 1'b0;  wr_cycle[  105] = 1'b1;  addr_rom[  105]='h000001a4;  wr_data_rom[  105]='h00000281;
    rd_cycle[  106] = 1'b0;  wr_cycle[  106] = 1'b1;  addr_rom[  106]='h000001a8;  wr_data_rom[  106]='h00000481;
    rd_cycle[  107] = 1'b0;  wr_cycle[  107] = 1'b1;  addr_rom[  107]='h000001ac;  wr_data_rom[  107]='h00000704;
    rd_cycle[  108] = 1'b0;  wr_cycle[  108] = 1'b1;  addr_rom[  108]='h000001b0;  wr_data_rom[  108]='h000007aa;
    rd_cycle[  109] = 1'b0;  wr_cycle[  109] = 1'b1;  addr_rom[  109]='h000001b4;  wr_data_rom[  109]='h00000504;
    rd_cycle[  110] = 1'b0;  wr_cycle[  110] = 1'b1;  addr_rom[  110]='h000001b8;  wr_data_rom[  110]='h00000035;
    rd_cycle[  111] = 1'b0;  wr_cycle[  111] = 1'b1;  addr_rom[  111]='h000001bc;  wr_data_rom[  111]='h00000504;
    rd_cycle[  112] = 1'b0;  wr_cycle[  112] = 1'b1;  addr_rom[  112]='h000001c0;  wr_data_rom[  112]='h000006bb;
    rd_cycle[  113] = 1'b0;  wr_cycle[  113] = 1'b1;  addr_rom[  113]='h000001c4;  wr_data_rom[  113]='h0000026e;
    rd_cycle[  114] = 1'b0;  wr_cycle[  114] = 1'b1;  addr_rom[  114]='h000001c8;  wr_data_rom[  114]='h00000534;
    rd_cycle[  115] = 1'b0;  wr_cycle[  115] = 1'b1;  addr_rom[  115]='h000001cc;  wr_data_rom[  115]='h00000627;
    rd_cycle[  116] = 1'b0;  wr_cycle[  116] = 1'b1;  addr_rom[  116]='h000001d0;  wr_data_rom[  116]='h000004ad;
    rd_cycle[  117] = 1'b0;  wr_cycle[  117] = 1'b1;  addr_rom[  117]='h000001d4;  wr_data_rom[  117]='h0000010a;
    rd_cycle[  118] = 1'b0;  wr_cycle[  118] = 1'b1;  addr_rom[  118]='h000001d8;  wr_data_rom[  118]='h0000030f;
    rd_cycle[  119] = 1'b0;  wr_cycle[  119] = 1'b1;  addr_rom[  119]='h000001dc;  wr_data_rom[  119]='h0000007e;
    rd_cycle[  120] = 1'b0;  wr_cycle[  120] = 1'b1;  addr_rom[  120]='h000001e0;  wr_data_rom[  120]='h00000441;
    rd_cycle[  121] = 1'b0;  wr_cycle[  121] = 1'b1;  addr_rom[  121]='h000001e4;  wr_data_rom[  121]='h00000071;
    rd_cycle[  122] = 1'b0;  wr_cycle[  122] = 1'b1;  addr_rom[  122]='h000001e8;  wr_data_rom[  122]='h000001f7;
    rd_cycle[  123] = 1'b0;  wr_cycle[  123] = 1'b1;  addr_rom[  123]='h000001ec;  wr_data_rom[  123]='h0000047f;
    rd_cycle[  124] = 1'b0;  wr_cycle[  124] = 1'b1;  addr_rom[  124]='h000001f0;  wr_data_rom[  124]='h000004fb;
    rd_cycle[  125] = 1'b0;  wr_cycle[  125] = 1'b1;  addr_rom[  125]='h000001f4;  wr_data_rom[  125]='h00000323;
    rd_cycle[  126] = 1'b0;  wr_cycle[  126] = 1'b1;  addr_rom[  126]='h000001f8;  wr_data_rom[  126]='h00000693;
    rd_cycle[  127] = 1'b0;  wr_cycle[  127] = 1'b1;  addr_rom[  127]='h000001fc;  wr_data_rom[  127]='h000004ab;
    rd_cycle[  128] = 1'b0;  wr_cycle[  128] = 1'b1;  addr_rom[  128]='h00000200;  wr_data_rom[  128]='h000007df;
    rd_cycle[  129] = 1'b0;  wr_cycle[  129] = 1'b1;  addr_rom[  129]='h00000204;  wr_data_rom[  129]='h000003dd;
    rd_cycle[  130] = 1'b0;  wr_cycle[  130] = 1'b1;  addr_rom[  130]='h00000208;  wr_data_rom[  130]='h0000028e;
    rd_cycle[  131] = 1'b0;  wr_cycle[  131] = 1'b1;  addr_rom[  131]='h0000020c;  wr_data_rom[  131]='h0000045e;
    rd_cycle[  132] = 1'b0;  wr_cycle[  132] = 1'b1;  addr_rom[  132]='h00000210;  wr_data_rom[  132]='h00000632;
    rd_cycle[  133] = 1'b0;  wr_cycle[  133] = 1'b1;  addr_rom[  133]='h00000214;  wr_data_rom[  133]='h000001d5;
    rd_cycle[  134] = 1'b0;  wr_cycle[  134] = 1'b1;  addr_rom[  134]='h00000218;  wr_data_rom[  134]='h00000674;
    rd_cycle[  135] = 1'b0;  wr_cycle[  135] = 1'b1;  addr_rom[  135]='h0000021c;  wr_data_rom[  135]='h000001e6;
    rd_cycle[  136] = 1'b0;  wr_cycle[  136] = 1'b1;  addr_rom[  136]='h00000220;  wr_data_rom[  136]='h0000079f;
    rd_cycle[  137] = 1'b0;  wr_cycle[  137] = 1'b1;  addr_rom[  137]='h00000224;  wr_data_rom[  137]='h000006e5;
    rd_cycle[  138] = 1'b0;  wr_cycle[  138] = 1'b1;  addr_rom[  138]='h00000228;  wr_data_rom[  138]='h000002e1;
    rd_cycle[  139] = 1'b0;  wr_cycle[  139] = 1'b1;  addr_rom[  139]='h0000022c;  wr_data_rom[  139]='h00000530;
    rd_cycle[  140] = 1'b0;  wr_cycle[  140] = 1'b1;  addr_rom[  140]='h00000230;  wr_data_rom[  140]='h0000032e;
    rd_cycle[  141] = 1'b0;  wr_cycle[  141] = 1'b1;  addr_rom[  141]='h00000234;  wr_data_rom[  141]='h00000588;
    rd_cycle[  142] = 1'b0;  wr_cycle[  142] = 1'b1;  addr_rom[  142]='h00000238;  wr_data_rom[  142]='h0000007d;
    rd_cycle[  143] = 1'b0;  wr_cycle[  143] = 1'b1;  addr_rom[  143]='h0000023c;  wr_data_rom[  143]='h000000df;
    rd_cycle[  144] = 1'b0;  wr_cycle[  144] = 1'b1;  addr_rom[  144]='h00000240;  wr_data_rom[  144]='h0000061e;
    rd_cycle[  145] = 1'b0;  wr_cycle[  145] = 1'b1;  addr_rom[  145]='h00000244;  wr_data_rom[  145]='h00000218;
    rd_cycle[  146] = 1'b0;  wr_cycle[  146] = 1'b1;  addr_rom[  146]='h00000248;  wr_data_rom[  146]='h000004d4;
    rd_cycle[  147] = 1'b0;  wr_cycle[  147] = 1'b1;  addr_rom[  147]='h0000024c;  wr_data_rom[  147]='h000001a3;
    rd_cycle[  148] = 1'b0;  wr_cycle[  148] = 1'b1;  addr_rom[  148]='h00000250;  wr_data_rom[  148]='h00000035;
    rd_cycle[  149] = 1'b0;  wr_cycle[  149] = 1'b1;  addr_rom[  149]='h00000254;  wr_data_rom[  149]='h000004b5;
    rd_cycle[  150] = 1'b0;  wr_cycle[  150] = 1'b1;  addr_rom[  150]='h00000258;  wr_data_rom[  150]='h000006e7;
    rd_cycle[  151] = 1'b0;  wr_cycle[  151] = 1'b1;  addr_rom[  151]='h0000025c;  wr_data_rom[  151]='h00000083;
    rd_cycle[  152] = 1'b0;  wr_cycle[  152] = 1'b1;  addr_rom[  152]='h00000260;  wr_data_rom[  152]='h000004fd;
    rd_cycle[  153] = 1'b0;  wr_cycle[  153] = 1'b1;  addr_rom[  153]='h00000264;  wr_data_rom[  153]='h00000624;
    rd_cycle[  154] = 1'b0;  wr_cycle[  154] = 1'b1;  addr_rom[  154]='h00000268;  wr_data_rom[  154]='h00000112;
    rd_cycle[  155] = 1'b0;  wr_cycle[  155] = 1'b1;  addr_rom[  155]='h0000026c;  wr_data_rom[  155]='h00000483;
    rd_cycle[  156] = 1'b0;  wr_cycle[  156] = 1'b1;  addr_rom[  156]='h00000270;  wr_data_rom[  156]='h000003ab;
    rd_cycle[  157] = 1'b0;  wr_cycle[  157] = 1'b1;  addr_rom[  157]='h00000274;  wr_data_rom[  157]='h000001dd;
    rd_cycle[  158] = 1'b0;  wr_cycle[  158] = 1'b1;  addr_rom[  158]='h00000278;  wr_data_rom[  158]='h000004f4;
    rd_cycle[  159] = 1'b0;  wr_cycle[  159] = 1'b1;  addr_rom[  159]='h0000027c;  wr_data_rom[  159]='h000005b9;
    rd_cycle[  160] = 1'b0;  wr_cycle[  160] = 1'b1;  addr_rom[  160]='h00000280;  wr_data_rom[  160]='h000007e9;
    rd_cycle[  161] = 1'b0;  wr_cycle[  161] = 1'b1;  addr_rom[  161]='h00000284;  wr_data_rom[  161]='h000002ff;
    rd_cycle[  162] = 1'b0;  wr_cycle[  162] = 1'b1;  addr_rom[  162]='h00000288;  wr_data_rom[  162]='h00000736;
    rd_cycle[  163] = 1'b0;  wr_cycle[  163] = 1'b1;  addr_rom[  163]='h0000028c;  wr_data_rom[  163]='h000002d9;
    rd_cycle[  164] = 1'b0;  wr_cycle[  164] = 1'b1;  addr_rom[  164]='h00000290;  wr_data_rom[  164]='h00000740;
    rd_cycle[  165] = 1'b0;  wr_cycle[  165] = 1'b1;  addr_rom[  165]='h00000294;  wr_data_rom[  165]='h0000012a;
    rd_cycle[  166] = 1'b0;  wr_cycle[  166] = 1'b1;  addr_rom[  166]='h00000298;  wr_data_rom[  166]='h00000699;
    rd_cycle[  167] = 1'b0;  wr_cycle[  167] = 1'b1;  addr_rom[  167]='h0000029c;  wr_data_rom[  167]='h0000073d;
    rd_cycle[  168] = 1'b0;  wr_cycle[  168] = 1'b1;  addr_rom[  168]='h000002a0;  wr_data_rom[  168]='h0000020d;
    rd_cycle[  169] = 1'b0;  wr_cycle[  169] = 1'b1;  addr_rom[  169]='h000002a4;  wr_data_rom[  169]='h0000014e;
    rd_cycle[  170] = 1'b0;  wr_cycle[  170] = 1'b1;  addr_rom[  170]='h000002a8;  wr_data_rom[  170]='h0000038a;
    rd_cycle[  171] = 1'b0;  wr_cycle[  171] = 1'b1;  addr_rom[  171]='h000002ac;  wr_data_rom[  171]='h00000376;
    rd_cycle[  172] = 1'b0;  wr_cycle[  172] = 1'b1;  addr_rom[  172]='h000002b0;  wr_data_rom[  172]='h00000380;
    rd_cycle[  173] = 1'b0;  wr_cycle[  173] = 1'b1;  addr_rom[  173]='h000002b4;  wr_data_rom[  173]='h00000288;
    rd_cycle[  174] = 1'b0;  wr_cycle[  174] = 1'b1;  addr_rom[  174]='h000002b8;  wr_data_rom[  174]='h00000479;
    rd_cycle[  175] = 1'b0;  wr_cycle[  175] = 1'b1;  addr_rom[  175]='h000002bc;  wr_data_rom[  175]='h00000542;
    rd_cycle[  176] = 1'b0;  wr_cycle[  176] = 1'b1;  addr_rom[  176]='h000002c0;  wr_data_rom[  176]='h000006c6;
    rd_cycle[  177] = 1'b0;  wr_cycle[  177] = 1'b1;  addr_rom[  177]='h000002c4;  wr_data_rom[  177]='h00000574;
    rd_cycle[  178] = 1'b0;  wr_cycle[  178] = 1'b1;  addr_rom[  178]='h000002c8;  wr_data_rom[  178]='h0000030e;
    rd_cycle[  179] = 1'b0;  wr_cycle[  179] = 1'b1;  addr_rom[  179]='h000002cc;  wr_data_rom[  179]='h0000003b;
    rd_cycle[  180] = 1'b0;  wr_cycle[  180] = 1'b1;  addr_rom[  180]='h000002d0;  wr_data_rom[  180]='h00000794;
    rd_cycle[  181] = 1'b0;  wr_cycle[  181] = 1'b1;  addr_rom[  181]='h000002d4;  wr_data_rom[  181]='h000003ef;
    rd_cycle[  182] = 1'b0;  wr_cycle[  182] = 1'b1;  addr_rom[  182]='h000002d8;  wr_data_rom[  182]='h000003db;
    rd_cycle[  183] = 1'b0;  wr_cycle[  183] = 1'b1;  addr_rom[  183]='h000002dc;  wr_data_rom[  183]='h0000012a;
    rd_cycle[  184] = 1'b0;  wr_cycle[  184] = 1'b1;  addr_rom[  184]='h000002e0;  wr_data_rom[  184]='h00000797;
    rd_cycle[  185] = 1'b0;  wr_cycle[  185] = 1'b1;  addr_rom[  185]='h000002e4;  wr_data_rom[  185]='h000003a0;
    rd_cycle[  186] = 1'b0;  wr_cycle[  186] = 1'b1;  addr_rom[  186]='h000002e8;  wr_data_rom[  186]='h000000da;
    rd_cycle[  187] = 1'b0;  wr_cycle[  187] = 1'b1;  addr_rom[  187]='h000002ec;  wr_data_rom[  187]='h0000067c;
    rd_cycle[  188] = 1'b0;  wr_cycle[  188] = 1'b1;  addr_rom[  188]='h000002f0;  wr_data_rom[  188]='h0000018d;
    rd_cycle[  189] = 1'b0;  wr_cycle[  189] = 1'b1;  addr_rom[  189]='h000002f4;  wr_data_rom[  189]='h00000336;
    rd_cycle[  190] = 1'b0;  wr_cycle[  190] = 1'b1;  addr_rom[  190]='h000002f8;  wr_data_rom[  190]='h000004dc;
    rd_cycle[  191] = 1'b0;  wr_cycle[  191] = 1'b1;  addr_rom[  191]='h000002fc;  wr_data_rom[  191]='h0000051d;
    rd_cycle[  192] = 1'b0;  wr_cycle[  192] = 1'b1;  addr_rom[  192]='h00000300;  wr_data_rom[  192]='h000004b0;
    rd_cycle[  193] = 1'b0;  wr_cycle[  193] = 1'b1;  addr_rom[  193]='h00000304;  wr_data_rom[  193]='h0000068a;
    rd_cycle[  194] = 1'b0;  wr_cycle[  194] = 1'b1;  addr_rom[  194]='h00000308;  wr_data_rom[  194]='h0000076c;
    rd_cycle[  195] = 1'b0;  wr_cycle[  195] = 1'b1;  addr_rom[  195]='h0000030c;  wr_data_rom[  195]='h000004f5;
    rd_cycle[  196] = 1'b0;  wr_cycle[  196] = 1'b1;  addr_rom[  196]='h00000310;  wr_data_rom[  196]='h00000544;
    rd_cycle[  197] = 1'b0;  wr_cycle[  197] = 1'b1;  addr_rom[  197]='h00000314;  wr_data_rom[  197]='h00000778;
    rd_cycle[  198] = 1'b0;  wr_cycle[  198] = 1'b1;  addr_rom[  198]='h00000318;  wr_data_rom[  198]='h0000060d;
    rd_cycle[  199] = 1'b0;  wr_cycle[  199] = 1'b1;  addr_rom[  199]='h0000031c;  wr_data_rom[  199]='h00000104;
    rd_cycle[  200] = 1'b0;  wr_cycle[  200] = 1'b1;  addr_rom[  200]='h00000320;  wr_data_rom[  200]='h00000741;
    rd_cycle[  201] = 1'b0;  wr_cycle[  201] = 1'b1;  addr_rom[  201]='h00000324;  wr_data_rom[  201]='h00000606;
    rd_cycle[  202] = 1'b0;  wr_cycle[  202] = 1'b1;  addr_rom[  202]='h00000328;  wr_data_rom[  202]='h000005a6;
    rd_cycle[  203] = 1'b0;  wr_cycle[  203] = 1'b1;  addr_rom[  203]='h0000032c;  wr_data_rom[  203]='h000006f8;
    rd_cycle[  204] = 1'b0;  wr_cycle[  204] = 1'b1;  addr_rom[  204]='h00000330;  wr_data_rom[  204]='h00000542;
    rd_cycle[  205] = 1'b0;  wr_cycle[  205] = 1'b1;  addr_rom[  205]='h00000334;  wr_data_rom[  205]='h0000079f;
    rd_cycle[  206] = 1'b0;  wr_cycle[  206] = 1'b1;  addr_rom[  206]='h00000338;  wr_data_rom[  206]='h00000670;
    rd_cycle[  207] = 1'b0;  wr_cycle[  207] = 1'b1;  addr_rom[  207]='h0000033c;  wr_data_rom[  207]='h000001ea;
    rd_cycle[  208] = 1'b0;  wr_cycle[  208] = 1'b1;  addr_rom[  208]='h00000340;  wr_data_rom[  208]='h0000077a;
    rd_cycle[  209] = 1'b0;  wr_cycle[  209] = 1'b1;  addr_rom[  209]='h00000344;  wr_data_rom[  209]='h000003a5;
    rd_cycle[  210] = 1'b0;  wr_cycle[  210] = 1'b1;  addr_rom[  210]='h00000348;  wr_data_rom[  210]='h000002c3;
    rd_cycle[  211] = 1'b0;  wr_cycle[  211] = 1'b1;  addr_rom[  211]='h0000034c;  wr_data_rom[  211]='h00000356;
    rd_cycle[  212] = 1'b0;  wr_cycle[  212] = 1'b1;  addr_rom[  212]='h00000350;  wr_data_rom[  212]='h000007ae;
    rd_cycle[  213] = 1'b0;  wr_cycle[  213] = 1'b1;  addr_rom[  213]='h00000354;  wr_data_rom[  213]='h00000116;
    rd_cycle[  214] = 1'b0;  wr_cycle[  214] = 1'b1;  addr_rom[  214]='h00000358;  wr_data_rom[  214]='h0000060c;
    rd_cycle[  215] = 1'b0;  wr_cycle[  215] = 1'b1;  addr_rom[  215]='h0000035c;  wr_data_rom[  215]='h000001f9;
    rd_cycle[  216] = 1'b0;  wr_cycle[  216] = 1'b1;  addr_rom[  216]='h00000360;  wr_data_rom[  216]='h00000120;
    rd_cycle[  217] = 1'b0;  wr_cycle[  217] = 1'b1;  addr_rom[  217]='h00000364;  wr_data_rom[  217]='h00000031;
    rd_cycle[  218] = 1'b0;  wr_cycle[  218] = 1'b1;  addr_rom[  218]='h00000368;  wr_data_rom[  218]='h000003bf;
    rd_cycle[  219] = 1'b0;  wr_cycle[  219] = 1'b1;  addr_rom[  219]='h0000036c;  wr_data_rom[  219]='h000006da;
    rd_cycle[  220] = 1'b0;  wr_cycle[  220] = 1'b1;  addr_rom[  220]='h00000370;  wr_data_rom[  220]='h0000046d;
    rd_cycle[  221] = 1'b0;  wr_cycle[  221] = 1'b1;  addr_rom[  221]='h00000374;  wr_data_rom[  221]='h00000338;
    rd_cycle[  222] = 1'b0;  wr_cycle[  222] = 1'b1;  addr_rom[  222]='h00000378;  wr_data_rom[  222]='h000000a5;
    rd_cycle[  223] = 1'b0;  wr_cycle[  223] = 1'b1;  addr_rom[  223]='h0000037c;  wr_data_rom[  223]='h00000568;
    rd_cycle[  224] = 1'b0;  wr_cycle[  224] = 1'b1;  addr_rom[  224]='h00000380;  wr_data_rom[  224]='h0000010f;
    rd_cycle[  225] = 1'b0;  wr_cycle[  225] = 1'b1;  addr_rom[  225]='h00000384;  wr_data_rom[  225]='h000006f9;
    rd_cycle[  226] = 1'b0;  wr_cycle[  226] = 1'b1;  addr_rom[  226]='h00000388;  wr_data_rom[  226]='h000006cb;
    rd_cycle[  227] = 1'b0;  wr_cycle[  227] = 1'b1;  addr_rom[  227]='h0000038c;  wr_data_rom[  227]='h00000747;
    rd_cycle[  228] = 1'b0;  wr_cycle[  228] = 1'b1;  addr_rom[  228]='h00000390;  wr_data_rom[  228]='h0000055e;
    rd_cycle[  229] = 1'b0;  wr_cycle[  229] = 1'b1;  addr_rom[  229]='h00000394;  wr_data_rom[  229]='h00000514;
    rd_cycle[  230] = 1'b0;  wr_cycle[  230] = 1'b1;  addr_rom[  230]='h00000398;  wr_data_rom[  230]='h000003d0;
    rd_cycle[  231] = 1'b0;  wr_cycle[  231] = 1'b1;  addr_rom[  231]='h0000039c;  wr_data_rom[  231]='h00000374;
    rd_cycle[  232] = 1'b0;  wr_cycle[  232] = 1'b1;  addr_rom[  232]='h000003a0;  wr_data_rom[  232]='h0000046a;
    rd_cycle[  233] = 1'b0;  wr_cycle[  233] = 1'b1;  addr_rom[  233]='h000003a4;  wr_data_rom[  233]='h000001a2;
    rd_cycle[  234] = 1'b0;  wr_cycle[  234] = 1'b1;  addr_rom[  234]='h000003a8;  wr_data_rom[  234]='h00000049;
    rd_cycle[  235] = 1'b0;  wr_cycle[  235] = 1'b1;  addr_rom[  235]='h000003ac;  wr_data_rom[  235]='h00000210;
    rd_cycle[  236] = 1'b0;  wr_cycle[  236] = 1'b1;  addr_rom[  236]='h000003b0;  wr_data_rom[  236]='h000004d0;
    rd_cycle[  237] = 1'b0;  wr_cycle[  237] = 1'b1;  addr_rom[  237]='h000003b4;  wr_data_rom[  237]='h0000078d;
    rd_cycle[  238] = 1'b0;  wr_cycle[  238] = 1'b1;  addr_rom[  238]='h000003b8;  wr_data_rom[  238]='h00000356;
    rd_cycle[  239] = 1'b0;  wr_cycle[  239] = 1'b1;  addr_rom[  239]='h000003bc;  wr_data_rom[  239]='h0000016c;
    rd_cycle[  240] = 1'b0;  wr_cycle[  240] = 1'b1;  addr_rom[  240]='h000003c0;  wr_data_rom[  240]='h000003a9;
    rd_cycle[  241] = 1'b0;  wr_cycle[  241] = 1'b1;  addr_rom[  241]='h000003c4;  wr_data_rom[  241]='h000000d6;
    rd_cycle[  242] = 1'b0;  wr_cycle[  242] = 1'b1;  addr_rom[  242]='h000003c8;  wr_data_rom[  242]='h0000028e;
    rd_cycle[  243] = 1'b0;  wr_cycle[  243] = 1'b1;  addr_rom[  243]='h000003cc;  wr_data_rom[  243]='h00000471;
    rd_cycle[  244] = 1'b0;  wr_cycle[  244] = 1'b1;  addr_rom[  244]='h000003d0;  wr_data_rom[  244]='h000005f2;
    rd_cycle[  245] = 1'b0;  wr_cycle[  245] = 1'b1;  addr_rom[  245]='h000003d4;  wr_data_rom[  245]='h0000001e;
    rd_cycle[  246] = 1'b0;  wr_cycle[  246] = 1'b1;  addr_rom[  246]='h000003d8;  wr_data_rom[  246]='h00000677;
    rd_cycle[  247] = 1'b0;  wr_cycle[  247] = 1'b1;  addr_rom[  247]='h000003dc;  wr_data_rom[  247]='h0000063f;
    rd_cycle[  248] = 1'b0;  wr_cycle[  248] = 1'b1;  addr_rom[  248]='h000003e0;  wr_data_rom[  248]='h000001df;
    rd_cycle[  249] = 1'b0;  wr_cycle[  249] = 1'b1;  addr_rom[  249]='h000003e4;  wr_data_rom[  249]='h000007d1;
    rd_cycle[  250] = 1'b0;  wr_cycle[  250] = 1'b1;  addr_rom[  250]='h000003e8;  wr_data_rom[  250]='h00000264;
    rd_cycle[  251] = 1'b0;  wr_cycle[  251] = 1'b1;  addr_rom[  251]='h000003ec;  wr_data_rom[  251]='h00000018;
    rd_cycle[  252] = 1'b0;  wr_cycle[  252] = 1'b1;  addr_rom[  252]='h000003f0;  wr_data_rom[  252]='h0000011f;
    rd_cycle[  253] = 1'b0;  wr_cycle[  253] = 1'b1;  addr_rom[  253]='h000003f4;  wr_data_rom[  253]='h0000005a;
    rd_cycle[  254] = 1'b0;  wr_cycle[  254] = 1'b1;  addr_rom[  254]='h000003f8;  wr_data_rom[  254]='h000004dd;
    rd_cycle[  255] = 1'b0;  wr_cycle[  255] = 1'b1;  addr_rom[  255]='h000003fc;  wr_data_rom[  255]='h0000064d;
    rd_cycle[  256] = 1'b0;  wr_cycle[  256] = 1'b1;  addr_rom[  256]='h00000400;  wr_data_rom[  256]='h00000379;
    rd_cycle[  257] = 1'b0;  wr_cycle[  257] = 1'b1;  addr_rom[  257]='h00000404;  wr_data_rom[  257]='h00000453;
    rd_cycle[  258] = 1'b0;  wr_cycle[  258] = 1'b1;  addr_rom[  258]='h00000408;  wr_data_rom[  258]='h00000288;
    rd_cycle[  259] = 1'b0;  wr_cycle[  259] = 1'b1;  addr_rom[  259]='h0000040c;  wr_data_rom[  259]='h000007d8;
    rd_cycle[  260] = 1'b0;  wr_cycle[  260] = 1'b1;  addr_rom[  260]='h00000410;  wr_data_rom[  260]='h000001a2;
    rd_cycle[  261] = 1'b0;  wr_cycle[  261] = 1'b1;  addr_rom[  261]='h00000414;  wr_data_rom[  261]='h000005e3;
    rd_cycle[  262] = 1'b0;  wr_cycle[  262] = 1'b1;  addr_rom[  262]='h00000418;  wr_data_rom[  262]='h00000513;
    rd_cycle[  263] = 1'b0;  wr_cycle[  263] = 1'b1;  addr_rom[  263]='h0000041c;  wr_data_rom[  263]='h0000054f;
    rd_cycle[  264] = 1'b0;  wr_cycle[  264] = 1'b1;  addr_rom[  264]='h00000420;  wr_data_rom[  264]='h000004ea;
    rd_cycle[  265] = 1'b0;  wr_cycle[  265] = 1'b1;  addr_rom[  265]='h00000424;  wr_data_rom[  265]='h000000bb;
    rd_cycle[  266] = 1'b0;  wr_cycle[  266] = 1'b1;  addr_rom[  266]='h00000428;  wr_data_rom[  266]='h0000029a;
    rd_cycle[  267] = 1'b0;  wr_cycle[  267] = 1'b1;  addr_rom[  267]='h0000042c;  wr_data_rom[  267]='h000005c2;
    rd_cycle[  268] = 1'b0;  wr_cycle[  268] = 1'b1;  addr_rom[  268]='h00000430;  wr_data_rom[  268]='h00000788;
    rd_cycle[  269] = 1'b0;  wr_cycle[  269] = 1'b1;  addr_rom[  269]='h00000434;  wr_data_rom[  269]='h000004a4;
    rd_cycle[  270] = 1'b0;  wr_cycle[  270] = 1'b1;  addr_rom[  270]='h00000438;  wr_data_rom[  270]='h000006cf;
    rd_cycle[  271] = 1'b0;  wr_cycle[  271] = 1'b1;  addr_rom[  271]='h0000043c;  wr_data_rom[  271]='h00000696;
    rd_cycle[  272] = 1'b0;  wr_cycle[  272] = 1'b1;  addr_rom[  272]='h00000440;  wr_data_rom[  272]='h00000410;
    rd_cycle[  273] = 1'b0;  wr_cycle[  273] = 1'b1;  addr_rom[  273]='h00000444;  wr_data_rom[  273]='h00000346;
    rd_cycle[  274] = 1'b0;  wr_cycle[  274] = 1'b1;  addr_rom[  274]='h00000448;  wr_data_rom[  274]='h00000282;
    rd_cycle[  275] = 1'b0;  wr_cycle[  275] = 1'b1;  addr_rom[  275]='h0000044c;  wr_data_rom[  275]='h000005dc;
    rd_cycle[  276] = 1'b0;  wr_cycle[  276] = 1'b1;  addr_rom[  276]='h00000450;  wr_data_rom[  276]='h000005fe;
    rd_cycle[  277] = 1'b0;  wr_cycle[  277] = 1'b1;  addr_rom[  277]='h00000454;  wr_data_rom[  277]='h00000273;
    rd_cycle[  278] = 1'b0;  wr_cycle[  278] = 1'b1;  addr_rom[  278]='h00000458;  wr_data_rom[  278]='h0000035c;
    rd_cycle[  279] = 1'b0;  wr_cycle[  279] = 1'b1;  addr_rom[  279]='h0000045c;  wr_data_rom[  279]='h000002c7;
    rd_cycle[  280] = 1'b0;  wr_cycle[  280] = 1'b1;  addr_rom[  280]='h00000460;  wr_data_rom[  280]='h00000228;
    rd_cycle[  281] = 1'b0;  wr_cycle[  281] = 1'b1;  addr_rom[  281]='h00000464;  wr_data_rom[  281]='h000003fc;
    rd_cycle[  282] = 1'b0;  wr_cycle[  282] = 1'b1;  addr_rom[  282]='h00000468;  wr_data_rom[  282]='h0000062c;
    rd_cycle[  283] = 1'b0;  wr_cycle[  283] = 1'b1;  addr_rom[  283]='h0000046c;  wr_data_rom[  283]='h00000605;
    rd_cycle[  284] = 1'b0;  wr_cycle[  284] = 1'b1;  addr_rom[  284]='h00000470;  wr_data_rom[  284]='h000004c4;
    rd_cycle[  285] = 1'b0;  wr_cycle[  285] = 1'b1;  addr_rom[  285]='h00000474;  wr_data_rom[  285]='h00000744;
    rd_cycle[  286] = 1'b0;  wr_cycle[  286] = 1'b1;  addr_rom[  286]='h00000478;  wr_data_rom[  286]='h0000034c;
    rd_cycle[  287] = 1'b0;  wr_cycle[  287] = 1'b1;  addr_rom[  287]='h0000047c;  wr_data_rom[  287]='h00000034;
    rd_cycle[  288] = 1'b0;  wr_cycle[  288] = 1'b1;  addr_rom[  288]='h00000480;  wr_data_rom[  288]='h0000026e;
    rd_cycle[  289] = 1'b0;  wr_cycle[  289] = 1'b1;  addr_rom[  289]='h00000484;  wr_data_rom[  289]='h000004ae;
    rd_cycle[  290] = 1'b0;  wr_cycle[  290] = 1'b1;  addr_rom[  290]='h00000488;  wr_data_rom[  290]='h000006fa;
    rd_cycle[  291] = 1'b0;  wr_cycle[  291] = 1'b1;  addr_rom[  291]='h0000048c;  wr_data_rom[  291]='h00000128;
    rd_cycle[  292] = 1'b0;  wr_cycle[  292] = 1'b1;  addr_rom[  292]='h00000490;  wr_data_rom[  292]='h00000143;
    rd_cycle[  293] = 1'b0;  wr_cycle[  293] = 1'b1;  addr_rom[  293]='h00000494;  wr_data_rom[  293]='h00000094;
    rd_cycle[  294] = 1'b0;  wr_cycle[  294] = 1'b1;  addr_rom[  294]='h00000498;  wr_data_rom[  294]='h000007b3;
    rd_cycle[  295] = 1'b0;  wr_cycle[  295] = 1'b1;  addr_rom[  295]='h0000049c;  wr_data_rom[  295]='h000007ca;
    rd_cycle[  296] = 1'b0;  wr_cycle[  296] = 1'b1;  addr_rom[  296]='h000004a0;  wr_data_rom[  296]='h0000055b;
    rd_cycle[  297] = 1'b0;  wr_cycle[  297] = 1'b1;  addr_rom[  297]='h000004a4;  wr_data_rom[  297]='h000006ea;
    rd_cycle[  298] = 1'b0;  wr_cycle[  298] = 1'b1;  addr_rom[  298]='h000004a8;  wr_data_rom[  298]='h000001bd;
    rd_cycle[  299] = 1'b0;  wr_cycle[  299] = 1'b1;  addr_rom[  299]='h000004ac;  wr_data_rom[  299]='h00000508;
    rd_cycle[  300] = 1'b0;  wr_cycle[  300] = 1'b1;  addr_rom[  300]='h000004b0;  wr_data_rom[  300]='h00000725;
    rd_cycle[  301] = 1'b0;  wr_cycle[  301] = 1'b1;  addr_rom[  301]='h000004b4;  wr_data_rom[  301]='h0000073a;
    rd_cycle[  302] = 1'b0;  wr_cycle[  302] = 1'b1;  addr_rom[  302]='h000004b8;  wr_data_rom[  302]='h0000026f;
    rd_cycle[  303] = 1'b0;  wr_cycle[  303] = 1'b1;  addr_rom[  303]='h000004bc;  wr_data_rom[  303]='h000002d7;
    rd_cycle[  304] = 1'b0;  wr_cycle[  304] = 1'b1;  addr_rom[  304]='h000004c0;  wr_data_rom[  304]='h0000004e;
    rd_cycle[  305] = 1'b0;  wr_cycle[  305] = 1'b1;  addr_rom[  305]='h000004c4;  wr_data_rom[  305]='h000002e3;
    rd_cycle[  306] = 1'b0;  wr_cycle[  306] = 1'b1;  addr_rom[  306]='h000004c8;  wr_data_rom[  306]='h00000235;
    rd_cycle[  307] = 1'b0;  wr_cycle[  307] = 1'b1;  addr_rom[  307]='h000004cc;  wr_data_rom[  307]='h00000302;
    rd_cycle[  308] = 1'b0;  wr_cycle[  308] = 1'b1;  addr_rom[  308]='h000004d0;  wr_data_rom[  308]='h00000706;
    rd_cycle[  309] = 1'b0;  wr_cycle[  309] = 1'b1;  addr_rom[  309]='h000004d4;  wr_data_rom[  309]='h0000001c;
    rd_cycle[  310] = 1'b0;  wr_cycle[  310] = 1'b1;  addr_rom[  310]='h000004d8;  wr_data_rom[  310]='h000006ba;
    rd_cycle[  311] = 1'b0;  wr_cycle[  311] = 1'b1;  addr_rom[  311]='h000004dc;  wr_data_rom[  311]='h00000313;
    rd_cycle[  312] = 1'b0;  wr_cycle[  312] = 1'b1;  addr_rom[  312]='h000004e0;  wr_data_rom[  312]='h00000712;
    rd_cycle[  313] = 1'b0;  wr_cycle[  313] = 1'b1;  addr_rom[  313]='h000004e4;  wr_data_rom[  313]='h00000618;
    rd_cycle[  314] = 1'b0;  wr_cycle[  314] = 1'b1;  addr_rom[  314]='h000004e8;  wr_data_rom[  314]='h00000619;
    rd_cycle[  315] = 1'b0;  wr_cycle[  315] = 1'b1;  addr_rom[  315]='h000004ec;  wr_data_rom[  315]='h000006a4;
    rd_cycle[  316] = 1'b0;  wr_cycle[  316] = 1'b1;  addr_rom[  316]='h000004f0;  wr_data_rom[  316]='h00000333;
    rd_cycle[  317] = 1'b0;  wr_cycle[  317] = 1'b1;  addr_rom[  317]='h000004f4;  wr_data_rom[  317]='h00000302;
    rd_cycle[  318] = 1'b0;  wr_cycle[  318] = 1'b1;  addr_rom[  318]='h000004f8;  wr_data_rom[  318]='h000005b1;
    rd_cycle[  319] = 1'b0;  wr_cycle[  319] = 1'b1;  addr_rom[  319]='h000004fc;  wr_data_rom[  319]='h00000755;
    rd_cycle[  320] = 1'b0;  wr_cycle[  320] = 1'b1;  addr_rom[  320]='h00000500;  wr_data_rom[  320]='h000005f9;
    rd_cycle[  321] = 1'b0;  wr_cycle[  321] = 1'b1;  addr_rom[  321]='h00000504;  wr_data_rom[  321]='h000005a3;
    rd_cycle[  322] = 1'b0;  wr_cycle[  322] = 1'b1;  addr_rom[  322]='h00000508;  wr_data_rom[  322]='h0000009c;
    rd_cycle[  323] = 1'b0;  wr_cycle[  323] = 1'b1;  addr_rom[  323]='h0000050c;  wr_data_rom[  323]='h00000726;
    rd_cycle[  324] = 1'b0;  wr_cycle[  324] = 1'b1;  addr_rom[  324]='h00000510;  wr_data_rom[  324]='h000007c5;
    rd_cycle[  325] = 1'b0;  wr_cycle[  325] = 1'b1;  addr_rom[  325]='h00000514;  wr_data_rom[  325]='h00000438;
    rd_cycle[  326] = 1'b0;  wr_cycle[  326] = 1'b1;  addr_rom[  326]='h00000518;  wr_data_rom[  326]='h0000009b;
    rd_cycle[  327] = 1'b0;  wr_cycle[  327] = 1'b1;  addr_rom[  327]='h0000051c;  wr_data_rom[  327]='h00000762;
    rd_cycle[  328] = 1'b0;  wr_cycle[  328] = 1'b1;  addr_rom[  328]='h00000520;  wr_data_rom[  328]='h00000221;
    rd_cycle[  329] = 1'b0;  wr_cycle[  329] = 1'b1;  addr_rom[  329]='h00000524;  wr_data_rom[  329]='h000000de;
    rd_cycle[  330] = 1'b0;  wr_cycle[  330] = 1'b1;  addr_rom[  330]='h00000528;  wr_data_rom[  330]='h000005c2;
    rd_cycle[  331] = 1'b0;  wr_cycle[  331] = 1'b1;  addr_rom[  331]='h0000052c;  wr_data_rom[  331]='h000006c7;
    rd_cycle[  332] = 1'b0;  wr_cycle[  332] = 1'b1;  addr_rom[  332]='h00000530;  wr_data_rom[  332]='h000003b1;
    rd_cycle[  333] = 1'b0;  wr_cycle[  333] = 1'b1;  addr_rom[  333]='h00000534;  wr_data_rom[  333]='h000005e6;
    rd_cycle[  334] = 1'b0;  wr_cycle[  334] = 1'b1;  addr_rom[  334]='h00000538;  wr_data_rom[  334]='h00000402;
    rd_cycle[  335] = 1'b0;  wr_cycle[  335] = 1'b1;  addr_rom[  335]='h0000053c;  wr_data_rom[  335]='h000003a3;
    rd_cycle[  336] = 1'b0;  wr_cycle[  336] = 1'b1;  addr_rom[  336]='h00000540;  wr_data_rom[  336]='h000000e5;
    rd_cycle[  337] = 1'b0;  wr_cycle[  337] = 1'b1;  addr_rom[  337]='h00000544;  wr_data_rom[  337]='h000002cb;
    rd_cycle[  338] = 1'b0;  wr_cycle[  338] = 1'b1;  addr_rom[  338]='h00000548;  wr_data_rom[  338]='h00000785;
    rd_cycle[  339] = 1'b0;  wr_cycle[  339] = 1'b1;  addr_rom[  339]='h0000054c;  wr_data_rom[  339]='h000002a1;
    rd_cycle[  340] = 1'b0;  wr_cycle[  340] = 1'b1;  addr_rom[  340]='h00000550;  wr_data_rom[  340]='h000005e5;
    rd_cycle[  341] = 1'b0;  wr_cycle[  341] = 1'b1;  addr_rom[  341]='h00000554;  wr_data_rom[  341]='h00000032;
    rd_cycle[  342] = 1'b0;  wr_cycle[  342] = 1'b1;  addr_rom[  342]='h00000558;  wr_data_rom[  342]='h000003d2;
    rd_cycle[  343] = 1'b0;  wr_cycle[  343] = 1'b1;  addr_rom[  343]='h0000055c;  wr_data_rom[  343]='h000006ab;
    rd_cycle[  344] = 1'b0;  wr_cycle[  344] = 1'b1;  addr_rom[  344]='h00000560;  wr_data_rom[  344]='h000000df;
    rd_cycle[  345] = 1'b0;  wr_cycle[  345] = 1'b1;  addr_rom[  345]='h00000564;  wr_data_rom[  345]='h000003f2;
    rd_cycle[  346] = 1'b0;  wr_cycle[  346] = 1'b1;  addr_rom[  346]='h00000568;  wr_data_rom[  346]='h00000124;
    rd_cycle[  347] = 1'b0;  wr_cycle[  347] = 1'b1;  addr_rom[  347]='h0000056c;  wr_data_rom[  347]='h000003fd;
    rd_cycle[  348] = 1'b0;  wr_cycle[  348] = 1'b1;  addr_rom[  348]='h00000570;  wr_data_rom[  348]='h00000432;
    rd_cycle[  349] = 1'b0;  wr_cycle[  349] = 1'b1;  addr_rom[  349]='h00000574;  wr_data_rom[  349]='h0000054e;
    rd_cycle[  350] = 1'b0;  wr_cycle[  350] = 1'b1;  addr_rom[  350]='h00000578;  wr_data_rom[  350]='h00000271;
    rd_cycle[  351] = 1'b0;  wr_cycle[  351] = 1'b1;  addr_rom[  351]='h0000057c;  wr_data_rom[  351]='h00000786;
    rd_cycle[  352] = 1'b0;  wr_cycle[  352] = 1'b1;  addr_rom[  352]='h00000580;  wr_data_rom[  352]='h00000103;
    rd_cycle[  353] = 1'b0;  wr_cycle[  353] = 1'b1;  addr_rom[  353]='h00000584;  wr_data_rom[  353]='h00000058;
    rd_cycle[  354] = 1'b0;  wr_cycle[  354] = 1'b1;  addr_rom[  354]='h00000588;  wr_data_rom[  354]='h00000122;
    rd_cycle[  355] = 1'b0;  wr_cycle[  355] = 1'b1;  addr_rom[  355]='h0000058c;  wr_data_rom[  355]='h000001b7;
    rd_cycle[  356] = 1'b0;  wr_cycle[  356] = 1'b1;  addr_rom[  356]='h00000590;  wr_data_rom[  356]='h00000543;
    rd_cycle[  357] = 1'b0;  wr_cycle[  357] = 1'b1;  addr_rom[  357]='h00000594;  wr_data_rom[  357]='h00000729;
    rd_cycle[  358] = 1'b0;  wr_cycle[  358] = 1'b1;  addr_rom[  358]='h00000598;  wr_data_rom[  358]='h00000351;
    rd_cycle[  359] = 1'b0;  wr_cycle[  359] = 1'b1;  addr_rom[  359]='h0000059c;  wr_data_rom[  359]='h000006ff;
    rd_cycle[  360] = 1'b0;  wr_cycle[  360] = 1'b1;  addr_rom[  360]='h000005a0;  wr_data_rom[  360]='h00000527;
    rd_cycle[  361] = 1'b0;  wr_cycle[  361] = 1'b1;  addr_rom[  361]='h000005a4;  wr_data_rom[  361]='h000007d2;
    rd_cycle[  362] = 1'b0;  wr_cycle[  362] = 1'b1;  addr_rom[  362]='h000005a8;  wr_data_rom[  362]='h00000149;
    rd_cycle[  363] = 1'b0;  wr_cycle[  363] = 1'b1;  addr_rom[  363]='h000005ac;  wr_data_rom[  363]='h00000225;
    rd_cycle[  364] = 1'b0;  wr_cycle[  364] = 1'b1;  addr_rom[  364]='h000005b0;  wr_data_rom[  364]='h00000642;
    rd_cycle[  365] = 1'b0;  wr_cycle[  365] = 1'b1;  addr_rom[  365]='h000005b4;  wr_data_rom[  365]='h00000266;
    rd_cycle[  366] = 1'b0;  wr_cycle[  366] = 1'b1;  addr_rom[  366]='h000005b8;  wr_data_rom[  366]='h000006d0;
    rd_cycle[  367] = 1'b0;  wr_cycle[  367] = 1'b1;  addr_rom[  367]='h000005bc;  wr_data_rom[  367]='h000003ac;
    rd_cycle[  368] = 1'b0;  wr_cycle[  368] = 1'b1;  addr_rom[  368]='h000005c0;  wr_data_rom[  368]='h0000031e;
    rd_cycle[  369] = 1'b0;  wr_cycle[  369] = 1'b1;  addr_rom[  369]='h000005c4;  wr_data_rom[  369]='h000000b7;
    rd_cycle[  370] = 1'b0;  wr_cycle[  370] = 1'b1;  addr_rom[  370]='h000005c8;  wr_data_rom[  370]='h0000042e;
    rd_cycle[  371] = 1'b0;  wr_cycle[  371] = 1'b1;  addr_rom[  371]='h000005cc;  wr_data_rom[  371]='h00000721;
    rd_cycle[  372] = 1'b0;  wr_cycle[  372] = 1'b1;  addr_rom[  372]='h000005d0;  wr_data_rom[  372]='h0000014b;
    rd_cycle[  373] = 1'b0;  wr_cycle[  373] = 1'b1;  addr_rom[  373]='h000005d4;  wr_data_rom[  373]='h00000434;
    rd_cycle[  374] = 1'b0;  wr_cycle[  374] = 1'b1;  addr_rom[  374]='h000005d8;  wr_data_rom[  374]='h0000078e;
    rd_cycle[  375] = 1'b0;  wr_cycle[  375] = 1'b1;  addr_rom[  375]='h000005dc;  wr_data_rom[  375]='h00000369;
    rd_cycle[  376] = 1'b0;  wr_cycle[  376] = 1'b1;  addr_rom[  376]='h000005e0;  wr_data_rom[  376]='h00000598;
    rd_cycle[  377] = 1'b0;  wr_cycle[  377] = 1'b1;  addr_rom[  377]='h000005e4;  wr_data_rom[  377]='h00000736;
    rd_cycle[  378] = 1'b0;  wr_cycle[  378] = 1'b1;  addr_rom[  378]='h000005e8;  wr_data_rom[  378]='h000007a1;
    rd_cycle[  379] = 1'b0;  wr_cycle[  379] = 1'b1;  addr_rom[  379]='h000005ec;  wr_data_rom[  379]='h00000439;
    rd_cycle[  380] = 1'b0;  wr_cycle[  380] = 1'b1;  addr_rom[  380]='h000005f0;  wr_data_rom[  380]='h000003f2;
    rd_cycle[  381] = 1'b0;  wr_cycle[  381] = 1'b1;  addr_rom[  381]='h000005f4;  wr_data_rom[  381]='h00000201;
    rd_cycle[  382] = 1'b0;  wr_cycle[  382] = 1'b1;  addr_rom[  382]='h000005f8;  wr_data_rom[  382]='h000002e7;
    rd_cycle[  383] = 1'b0;  wr_cycle[  383] = 1'b1;  addr_rom[  383]='h000005fc;  wr_data_rom[  383]='h000002a1;
    rd_cycle[  384] = 1'b0;  wr_cycle[  384] = 1'b1;  addr_rom[  384]='h00000600;  wr_data_rom[  384]='h0000001c;
    rd_cycle[  385] = 1'b0;  wr_cycle[  385] = 1'b1;  addr_rom[  385]='h00000604;  wr_data_rom[  385]='h0000056c;
    rd_cycle[  386] = 1'b0;  wr_cycle[  386] = 1'b1;  addr_rom[  386]='h00000608;  wr_data_rom[  386]='h0000011a;
    rd_cycle[  387] = 1'b0;  wr_cycle[  387] = 1'b1;  addr_rom[  387]='h0000060c;  wr_data_rom[  387]='h000004c6;
    rd_cycle[  388] = 1'b0;  wr_cycle[  388] = 1'b1;  addr_rom[  388]='h00000610;  wr_data_rom[  388]='h000002ad;
    rd_cycle[  389] = 1'b0;  wr_cycle[  389] = 1'b1;  addr_rom[  389]='h00000614;  wr_data_rom[  389]='h0000067a;
    rd_cycle[  390] = 1'b0;  wr_cycle[  390] = 1'b1;  addr_rom[  390]='h00000618;  wr_data_rom[  390]='h000004a9;
    rd_cycle[  391] = 1'b0;  wr_cycle[  391] = 1'b1;  addr_rom[  391]='h0000061c;  wr_data_rom[  391]='h00000355;
    rd_cycle[  392] = 1'b0;  wr_cycle[  392] = 1'b1;  addr_rom[  392]='h00000620;  wr_data_rom[  392]='h0000069b;
    rd_cycle[  393] = 1'b0;  wr_cycle[  393] = 1'b1;  addr_rom[  393]='h00000624;  wr_data_rom[  393]='h000007a4;
    rd_cycle[  394] = 1'b0;  wr_cycle[  394] = 1'b1;  addr_rom[  394]='h00000628;  wr_data_rom[  394]='h00000294;
    rd_cycle[  395] = 1'b0;  wr_cycle[  395] = 1'b1;  addr_rom[  395]='h0000062c;  wr_data_rom[  395]='h0000009c;
    rd_cycle[  396] = 1'b0;  wr_cycle[  396] = 1'b1;  addr_rom[  396]='h00000630;  wr_data_rom[  396]='h00000526;
    rd_cycle[  397] = 1'b0;  wr_cycle[  397] = 1'b1;  addr_rom[  397]='h00000634;  wr_data_rom[  397]='h000000f1;
    rd_cycle[  398] = 1'b0;  wr_cycle[  398] = 1'b1;  addr_rom[  398]='h00000638;  wr_data_rom[  398]='h00000161;
    rd_cycle[  399] = 1'b0;  wr_cycle[  399] = 1'b1;  addr_rom[  399]='h0000063c;  wr_data_rom[  399]='h000007e9;
    rd_cycle[  400] = 1'b0;  wr_cycle[  400] = 1'b1;  addr_rom[  400]='h00000640;  wr_data_rom[  400]='h00000048;
    rd_cycle[  401] = 1'b0;  wr_cycle[  401] = 1'b1;  addr_rom[  401]='h00000644;  wr_data_rom[  401]='h000004a0;
    rd_cycle[  402] = 1'b0;  wr_cycle[  402] = 1'b1;  addr_rom[  402]='h00000648;  wr_data_rom[  402]='h0000029c;
    rd_cycle[  403] = 1'b0;  wr_cycle[  403] = 1'b1;  addr_rom[  403]='h0000064c;  wr_data_rom[  403]='h000006a2;
    rd_cycle[  404] = 1'b0;  wr_cycle[  404] = 1'b1;  addr_rom[  404]='h00000650;  wr_data_rom[  404]='h000003ff;
    rd_cycle[  405] = 1'b0;  wr_cycle[  405] = 1'b1;  addr_rom[  405]='h00000654;  wr_data_rom[  405]='h0000045f;
    rd_cycle[  406] = 1'b0;  wr_cycle[  406] = 1'b1;  addr_rom[  406]='h00000658;  wr_data_rom[  406]='h00000669;
    rd_cycle[  407] = 1'b0;  wr_cycle[  407] = 1'b1;  addr_rom[  407]='h0000065c;  wr_data_rom[  407]='h000005cc;
    rd_cycle[  408] = 1'b0;  wr_cycle[  408] = 1'b1;  addr_rom[  408]='h00000660;  wr_data_rom[  408]='h0000077c;
    rd_cycle[  409] = 1'b0;  wr_cycle[  409] = 1'b1;  addr_rom[  409]='h00000664;  wr_data_rom[  409]='h000006f8;
    rd_cycle[  410] = 1'b0;  wr_cycle[  410] = 1'b1;  addr_rom[  410]='h00000668;  wr_data_rom[  410]='h000007cf;
    rd_cycle[  411] = 1'b0;  wr_cycle[  411] = 1'b1;  addr_rom[  411]='h0000066c;  wr_data_rom[  411]='h0000017e;
    rd_cycle[  412] = 1'b0;  wr_cycle[  412] = 1'b1;  addr_rom[  412]='h00000670;  wr_data_rom[  412]='h000000a8;
    rd_cycle[  413] = 1'b0;  wr_cycle[  413] = 1'b1;  addr_rom[  413]='h00000674;  wr_data_rom[  413]='h00000354;
    rd_cycle[  414] = 1'b0;  wr_cycle[  414] = 1'b1;  addr_rom[  414]='h00000678;  wr_data_rom[  414]='h000007ea;
    rd_cycle[  415] = 1'b0;  wr_cycle[  415] = 1'b1;  addr_rom[  415]='h0000067c;  wr_data_rom[  415]='h00000274;
    rd_cycle[  416] = 1'b0;  wr_cycle[  416] = 1'b1;  addr_rom[  416]='h00000680;  wr_data_rom[  416]='h000002f5;
    rd_cycle[  417] = 1'b0;  wr_cycle[  417] = 1'b1;  addr_rom[  417]='h00000684;  wr_data_rom[  417]='h0000073c;
    rd_cycle[  418] = 1'b0;  wr_cycle[  418] = 1'b1;  addr_rom[  418]='h00000688;  wr_data_rom[  418]='h0000054a;
    rd_cycle[  419] = 1'b0;  wr_cycle[  419] = 1'b1;  addr_rom[  419]='h0000068c;  wr_data_rom[  419]='h0000040c;
    rd_cycle[  420] = 1'b0;  wr_cycle[  420] = 1'b1;  addr_rom[  420]='h00000690;  wr_data_rom[  420]='h00000554;
    rd_cycle[  421] = 1'b0;  wr_cycle[  421] = 1'b1;  addr_rom[  421]='h00000694;  wr_data_rom[  421]='h00000506;
    rd_cycle[  422] = 1'b0;  wr_cycle[  422] = 1'b1;  addr_rom[  422]='h00000698;  wr_data_rom[  422]='h000002d9;
    rd_cycle[  423] = 1'b0;  wr_cycle[  423] = 1'b1;  addr_rom[  423]='h0000069c;  wr_data_rom[  423]='h000004a7;
    rd_cycle[  424] = 1'b0;  wr_cycle[  424] = 1'b1;  addr_rom[  424]='h000006a0;  wr_data_rom[  424]='h0000037a;
    rd_cycle[  425] = 1'b0;  wr_cycle[  425] = 1'b1;  addr_rom[  425]='h000006a4;  wr_data_rom[  425]='h00000153;
    rd_cycle[  426] = 1'b0;  wr_cycle[  426] = 1'b1;  addr_rom[  426]='h000006a8;  wr_data_rom[  426]='h00000136;
    rd_cycle[  427] = 1'b0;  wr_cycle[  427] = 1'b1;  addr_rom[  427]='h000006ac;  wr_data_rom[  427]='h000001ab;
    rd_cycle[  428] = 1'b0;  wr_cycle[  428] = 1'b1;  addr_rom[  428]='h000006b0;  wr_data_rom[  428]='h0000056e;
    rd_cycle[  429] = 1'b0;  wr_cycle[  429] = 1'b1;  addr_rom[  429]='h000006b4;  wr_data_rom[  429]='h0000034b;
    rd_cycle[  430] = 1'b0;  wr_cycle[  430] = 1'b1;  addr_rom[  430]='h000006b8;  wr_data_rom[  430]='h000007ad;
    rd_cycle[  431] = 1'b0;  wr_cycle[  431] = 1'b1;  addr_rom[  431]='h000006bc;  wr_data_rom[  431]='h000001ef;
    rd_cycle[  432] = 1'b0;  wr_cycle[  432] = 1'b1;  addr_rom[  432]='h000006c0;  wr_data_rom[  432]='h00000654;
    rd_cycle[  433] = 1'b0;  wr_cycle[  433] = 1'b1;  addr_rom[  433]='h000006c4;  wr_data_rom[  433]='h00000314;
    rd_cycle[  434] = 1'b0;  wr_cycle[  434] = 1'b1;  addr_rom[  434]='h000006c8;  wr_data_rom[  434]='h000000f3;
    rd_cycle[  435] = 1'b0;  wr_cycle[  435] = 1'b1;  addr_rom[  435]='h000006cc;  wr_data_rom[  435]='h0000011e;
    rd_cycle[  436] = 1'b0;  wr_cycle[  436] = 1'b1;  addr_rom[  436]='h000006d0;  wr_data_rom[  436]='h0000037d;
    rd_cycle[  437] = 1'b0;  wr_cycle[  437] = 1'b1;  addr_rom[  437]='h000006d4;  wr_data_rom[  437]='h000000f6;
    rd_cycle[  438] = 1'b0;  wr_cycle[  438] = 1'b1;  addr_rom[  438]='h000006d8;  wr_data_rom[  438]='h00000059;
    rd_cycle[  439] = 1'b0;  wr_cycle[  439] = 1'b1;  addr_rom[  439]='h000006dc;  wr_data_rom[  439]='h0000055f;
    rd_cycle[  440] = 1'b0;  wr_cycle[  440] = 1'b1;  addr_rom[  440]='h000006e0;  wr_data_rom[  440]='h000006c8;
    rd_cycle[  441] = 1'b0;  wr_cycle[  441] = 1'b1;  addr_rom[  441]='h000006e4;  wr_data_rom[  441]='h0000010e;
    rd_cycle[  442] = 1'b0;  wr_cycle[  442] = 1'b1;  addr_rom[  442]='h000006e8;  wr_data_rom[  442]='h000000a1;
    rd_cycle[  443] = 1'b0;  wr_cycle[  443] = 1'b1;  addr_rom[  443]='h000006ec;  wr_data_rom[  443]='h0000057b;
    rd_cycle[  444] = 1'b0;  wr_cycle[  444] = 1'b1;  addr_rom[  444]='h000006f0;  wr_data_rom[  444]='h00000146;
    rd_cycle[  445] = 1'b0;  wr_cycle[  445] = 1'b1;  addr_rom[  445]='h000006f4;  wr_data_rom[  445]='h000003ca;
    rd_cycle[  446] = 1'b0;  wr_cycle[  446] = 1'b1;  addr_rom[  446]='h000006f8;  wr_data_rom[  446]='h00000150;
    rd_cycle[  447] = 1'b0;  wr_cycle[  447] = 1'b1;  addr_rom[  447]='h000006fc;  wr_data_rom[  447]='h000002a7;
    rd_cycle[  448] = 1'b0;  wr_cycle[  448] = 1'b1;  addr_rom[  448]='h00000700;  wr_data_rom[  448]='h00000225;
    rd_cycle[  449] = 1'b0;  wr_cycle[  449] = 1'b1;  addr_rom[  449]='h00000704;  wr_data_rom[  449]='h000003b2;
    rd_cycle[  450] = 1'b0;  wr_cycle[  450] = 1'b1;  addr_rom[  450]='h00000708;  wr_data_rom[  450]='h00000125;
    rd_cycle[  451] = 1'b0;  wr_cycle[  451] = 1'b1;  addr_rom[  451]='h0000070c;  wr_data_rom[  451]='h000006c8;
    rd_cycle[  452] = 1'b0;  wr_cycle[  452] = 1'b1;  addr_rom[  452]='h00000710;  wr_data_rom[  452]='h0000074f;
    rd_cycle[  453] = 1'b0;  wr_cycle[  453] = 1'b1;  addr_rom[  453]='h00000714;  wr_data_rom[  453]='h000002ac;
    rd_cycle[  454] = 1'b0;  wr_cycle[  454] = 1'b1;  addr_rom[  454]='h00000718;  wr_data_rom[  454]='h000002e1;
    rd_cycle[  455] = 1'b0;  wr_cycle[  455] = 1'b1;  addr_rom[  455]='h0000071c;  wr_data_rom[  455]='h0000053b;
    rd_cycle[  456] = 1'b0;  wr_cycle[  456] = 1'b1;  addr_rom[  456]='h00000720;  wr_data_rom[  456]='h0000062c;
    rd_cycle[  457] = 1'b0;  wr_cycle[  457] = 1'b1;  addr_rom[  457]='h00000724;  wr_data_rom[  457]='h00000193;
    rd_cycle[  458] = 1'b0;  wr_cycle[  458] = 1'b1;  addr_rom[  458]='h00000728;  wr_data_rom[  458]='h0000028a;
    rd_cycle[  459] = 1'b0;  wr_cycle[  459] = 1'b1;  addr_rom[  459]='h0000072c;  wr_data_rom[  459]='h00000506;
    rd_cycle[  460] = 1'b0;  wr_cycle[  460] = 1'b1;  addr_rom[  460]='h00000730;  wr_data_rom[  460]='h00000005;
    rd_cycle[  461] = 1'b0;  wr_cycle[  461] = 1'b1;  addr_rom[  461]='h00000734;  wr_data_rom[  461]='h000007cd;
    rd_cycle[  462] = 1'b0;  wr_cycle[  462] = 1'b1;  addr_rom[  462]='h00000738;  wr_data_rom[  462]='h000000b9;
    rd_cycle[  463] = 1'b0;  wr_cycle[  463] = 1'b1;  addr_rom[  463]='h0000073c;  wr_data_rom[  463]='h000005fc;
    rd_cycle[  464] = 1'b0;  wr_cycle[  464] = 1'b1;  addr_rom[  464]='h00000740;  wr_data_rom[  464]='h000004db;
    rd_cycle[  465] = 1'b0;  wr_cycle[  465] = 1'b1;  addr_rom[  465]='h00000744;  wr_data_rom[  465]='h000004b2;
    rd_cycle[  466] = 1'b0;  wr_cycle[  466] = 1'b1;  addr_rom[  466]='h00000748;  wr_data_rom[  466]='h00000704;
    rd_cycle[  467] = 1'b0;  wr_cycle[  467] = 1'b1;  addr_rom[  467]='h0000074c;  wr_data_rom[  467]='h000004a5;
    rd_cycle[  468] = 1'b0;  wr_cycle[  468] = 1'b1;  addr_rom[  468]='h00000750;  wr_data_rom[  468]='h000004d5;
    rd_cycle[  469] = 1'b0;  wr_cycle[  469] = 1'b1;  addr_rom[  469]='h00000754;  wr_data_rom[  469]='h00000010;
    rd_cycle[  470] = 1'b0;  wr_cycle[  470] = 1'b1;  addr_rom[  470]='h00000758;  wr_data_rom[  470]='h00000721;
    rd_cycle[  471] = 1'b0;  wr_cycle[  471] = 1'b1;  addr_rom[  471]='h0000075c;  wr_data_rom[  471]='h000003fc;
    rd_cycle[  472] = 1'b0;  wr_cycle[  472] = 1'b1;  addr_rom[  472]='h00000760;  wr_data_rom[  472]='h00000398;
    rd_cycle[  473] = 1'b0;  wr_cycle[  473] = 1'b1;  addr_rom[  473]='h00000764;  wr_data_rom[  473]='h0000025f;
    rd_cycle[  474] = 1'b0;  wr_cycle[  474] = 1'b1;  addr_rom[  474]='h00000768;  wr_data_rom[  474]='h000002b0;
    rd_cycle[  475] = 1'b0;  wr_cycle[  475] = 1'b1;  addr_rom[  475]='h0000076c;  wr_data_rom[  475]='h000004a2;
    rd_cycle[  476] = 1'b0;  wr_cycle[  476] = 1'b1;  addr_rom[  476]='h00000770;  wr_data_rom[  476]='h0000003d;
    rd_cycle[  477] = 1'b0;  wr_cycle[  477] = 1'b1;  addr_rom[  477]='h00000774;  wr_data_rom[  477]='h0000018c;
    rd_cycle[  478] = 1'b0;  wr_cycle[  478] = 1'b1;  addr_rom[  478]='h00000778;  wr_data_rom[  478]='h00000525;
    rd_cycle[  479] = 1'b0;  wr_cycle[  479] = 1'b1;  addr_rom[  479]='h0000077c;  wr_data_rom[  479]='h000002b5;
    rd_cycle[  480] = 1'b0;  wr_cycle[  480] = 1'b1;  addr_rom[  480]='h00000780;  wr_data_rom[  480]='h00000330;
    rd_cycle[  481] = 1'b0;  wr_cycle[  481] = 1'b1;  addr_rom[  481]='h00000784;  wr_data_rom[  481]='h000004db;
    rd_cycle[  482] = 1'b0;  wr_cycle[  482] = 1'b1;  addr_rom[  482]='h00000788;  wr_data_rom[  482]='h00000574;
    rd_cycle[  483] = 1'b0;  wr_cycle[  483] = 1'b1;  addr_rom[  483]='h0000078c;  wr_data_rom[  483]='h000002bf;
    rd_cycle[  484] = 1'b0;  wr_cycle[  484] = 1'b1;  addr_rom[  484]='h00000790;  wr_data_rom[  484]='h000006d6;
    rd_cycle[  485] = 1'b0;  wr_cycle[  485] = 1'b1;  addr_rom[  485]='h00000794;  wr_data_rom[  485]='h0000044f;
    rd_cycle[  486] = 1'b0;  wr_cycle[  486] = 1'b1;  addr_rom[  486]='h00000798;  wr_data_rom[  486]='h00000131;
    rd_cycle[  487] = 1'b0;  wr_cycle[  487] = 1'b1;  addr_rom[  487]='h0000079c;  wr_data_rom[  487]='h0000039c;
    rd_cycle[  488] = 1'b0;  wr_cycle[  488] = 1'b1;  addr_rom[  488]='h000007a0;  wr_data_rom[  488]='h0000034f;
    rd_cycle[  489] = 1'b0;  wr_cycle[  489] = 1'b1;  addr_rom[  489]='h000007a4;  wr_data_rom[  489]='h000001e7;
    rd_cycle[  490] = 1'b0;  wr_cycle[  490] = 1'b1;  addr_rom[  490]='h000007a8;  wr_data_rom[  490]='h000003d9;
    rd_cycle[  491] = 1'b0;  wr_cycle[  491] = 1'b1;  addr_rom[  491]='h000007ac;  wr_data_rom[  491]='h0000021f;
    rd_cycle[  492] = 1'b0;  wr_cycle[  492] = 1'b1;  addr_rom[  492]='h000007b0;  wr_data_rom[  492]='h000003b0;
    rd_cycle[  493] = 1'b0;  wr_cycle[  493] = 1'b1;  addr_rom[  493]='h000007b4;  wr_data_rom[  493]='h00000576;
    rd_cycle[  494] = 1'b0;  wr_cycle[  494] = 1'b1;  addr_rom[  494]='h000007b8;  wr_data_rom[  494]='h000002ab;
    rd_cycle[  495] = 1'b0;  wr_cycle[  495] = 1'b1;  addr_rom[  495]='h000007bc;  wr_data_rom[  495]='h00000343;
    rd_cycle[  496] = 1'b0;  wr_cycle[  496] = 1'b1;  addr_rom[  496]='h000007c0;  wr_data_rom[  496]='h000002c4;
    rd_cycle[  497] = 1'b0;  wr_cycle[  497] = 1'b1;  addr_rom[  497]='h000007c4;  wr_data_rom[  497]='h0000024b;
    rd_cycle[  498] = 1'b0;  wr_cycle[  498] = 1'b1;  addr_rom[  498]='h000007c8;  wr_data_rom[  498]='h00000168;
    rd_cycle[  499] = 1'b0;  wr_cycle[  499] = 1'b1;  addr_rom[  499]='h000007cc;  wr_data_rom[  499]='h0000065c;
    rd_cycle[  500] = 1'b0;  wr_cycle[  500] = 1'b1;  addr_rom[  500]='h000007d0;  wr_data_rom[  500]='h000004aa;
    rd_cycle[  501] = 1'b0;  wr_cycle[  501] = 1'b1;  addr_rom[  501]='h000007d4;  wr_data_rom[  501]='h0000007d;
    rd_cycle[  502] = 1'b0;  wr_cycle[  502] = 1'b1;  addr_rom[  502]='h000007d8;  wr_data_rom[  502]='h0000028f;
    rd_cycle[  503] = 1'b0;  wr_cycle[  503] = 1'b1;  addr_rom[  503]='h000007dc;  wr_data_rom[  503]='h000005cb;
    rd_cycle[  504] = 1'b0;  wr_cycle[  504] = 1'b1;  addr_rom[  504]='h000007e0;  wr_data_rom[  504]='h0000052b;
    rd_cycle[  505] = 1'b0;  wr_cycle[  505] = 1'b1;  addr_rom[  505]='h000007e4;  wr_data_rom[  505]='h00000347;
    rd_cycle[  506] = 1'b0;  wr_cycle[  506] = 1'b1;  addr_rom[  506]='h000007e8;  wr_data_rom[  506]='h00000180;
    rd_cycle[  507] = 1'b0;  wr_cycle[  507] = 1'b1;  addr_rom[  507]='h000007ec;  wr_data_rom[  507]='h00000096;
    rd_cycle[  508] = 1'b0;  wr_cycle[  508] = 1'b1;  addr_rom[  508]='h000007f0;  wr_data_rom[  508]='h00000035;
    rd_cycle[  509] = 1'b0;  wr_cycle[  509] = 1'b1;  addr_rom[  509]='h000007f4;  wr_data_rom[  509]='h000005a9;
    rd_cycle[  510] = 1'b0;  wr_cycle[  510] = 1'b1;  addr_rom[  510]='h000007f8;  wr_data_rom[  510]='h00000400;
    rd_cycle[  511] = 1'b0;  wr_cycle[  511] = 1'b1;  addr_rom[  511]='h000007fc;  wr_data_rom[  511]='h000000fd;
    // 1536 random read and write cycles
    rd_cycle[  512] = 1'b1;  wr_cycle[  512] = 1'b0;  addr_rom[  512]='h000005f8;  wr_data_rom[  512]='h00000000;
    rd_cycle[  513] = 1'b1;  wr_cycle[  513] = 1'b0;  addr_rom[  513]='h000006c8;  wr_data_rom[  513]='h00000000;
    rd_cycle[  514] = 1'b0;  wr_cycle[  514] = 1'b1;  addr_rom[  514]='h000007c4;  wr_data_rom[  514]='h000000da;
    rd_cycle[  515] = 1'b0;  wr_cycle[  515] = 1'b1;  addr_rom[  515]='h00000128;  wr_data_rom[  515]='h00000007;
    rd_cycle[  516] = 1'b0;  wr_cycle[  516] = 1'b1;  addr_rom[  516]='h000005dc;  wr_data_rom[  516]='h00000480;
    rd_cycle[  517] = 1'b1;  wr_cycle[  517] = 1'b0;  addr_rom[  517]='h00000320;  wr_data_rom[  517]='h00000000;
    rd_cycle[  518] = 1'b1;  wr_cycle[  518] = 1'b0;  addr_rom[  518]='h00000130;  wr_data_rom[  518]='h00000000;
    rd_cycle[  519] = 1'b1;  wr_cycle[  519] = 1'b0;  addr_rom[  519]='h0000041c;  wr_data_rom[  519]='h00000000;
    rd_cycle[  520] = 1'b0;  wr_cycle[  520] = 1'b1;  addr_rom[  520]='h00000210;  wr_data_rom[  520]='h00000468;
    rd_cycle[  521] = 1'b1;  wr_cycle[  521] = 1'b0;  addr_rom[  521]='h000005b8;  wr_data_rom[  521]='h00000000;
    rd_cycle[  522] = 1'b0;  wr_cycle[  522] = 1'b1;  addr_rom[  522]='h000003b8;  wr_data_rom[  522]='h000001d6;
    rd_cycle[  523] = 1'b1;  wr_cycle[  523] = 1'b0;  addr_rom[  523]='h00000220;  wr_data_rom[  523]='h00000000;
    rd_cycle[  524] = 1'b0;  wr_cycle[  524] = 1'b1;  addr_rom[  524]='h00000034;  wr_data_rom[  524]='h000005ef;
    rd_cycle[  525] = 1'b0;  wr_cycle[  525] = 1'b1;  addr_rom[  525]='h00000024;  wr_data_rom[  525]='h00000646;
    rd_cycle[  526] = 1'b0;  wr_cycle[  526] = 1'b1;  addr_rom[  526]='h00000640;  wr_data_rom[  526]='h000007e7;
    rd_cycle[  527] = 1'b1;  wr_cycle[  527] = 1'b0;  addr_rom[  527]='h0000051c;  wr_data_rom[  527]='h00000000;
    rd_cycle[  528] = 1'b1;  wr_cycle[  528] = 1'b0;  addr_rom[  528]='h00000310;  wr_data_rom[  528]='h00000000;
    rd_cycle[  529] = 1'b0;  wr_cycle[  529] = 1'b1;  addr_rom[  529]='h000006d4;  wr_data_rom[  529]='h000000ce;
    rd_cycle[  530] = 1'b0;  wr_cycle[  530] = 1'b1;  addr_rom[  530]='h0000045c;  wr_data_rom[  530]='h000004f4;
    rd_cycle[  531] = 1'b0;  wr_cycle[  531] = 1'b1;  addr_rom[  531]='h000005c4;  wr_data_rom[  531]='h00000192;
    rd_cycle[  532] = 1'b0;  wr_cycle[  532] = 1'b1;  addr_rom[  532]='h00000108;  wr_data_rom[  532]='h000003b1;
    rd_cycle[  533] = 1'b0;  wr_cycle[  533] = 1'b1;  addr_rom[  533]='h000002c0;  wr_data_rom[  533]='h000004a9;
    rd_cycle[  534] = 1'b1;  wr_cycle[  534] = 1'b0;  addr_rom[  534]='h0000014c;  wr_data_rom[  534]='h00000000;
    rd_cycle[  535] = 1'b1;  wr_cycle[  535] = 1'b0;  addr_rom[  535]='h00000754;  wr_data_rom[  535]='h00000000;
    rd_cycle[  536] = 1'b1;  wr_cycle[  536] = 1'b0;  addr_rom[  536]='h0000073c;  wr_data_rom[  536]='h00000000;
    rd_cycle[  537] = 1'b0;  wr_cycle[  537] = 1'b1;  addr_rom[  537]='h000004ec;  wr_data_rom[  537]='h000005cb;
    rd_cycle[  538] = 1'b0;  wr_cycle[  538] = 1'b1;  addr_rom[  538]='h00000608;  wr_data_rom[  538]='h000004f2;
    rd_cycle[  539] = 1'b1;  wr_cycle[  539] = 1'b0;  addr_rom[  539]='h000000a4;  wr_data_rom[  539]='h00000000;
    rd_cycle[  540] = 1'b0;  wr_cycle[  540] = 1'b1;  addr_rom[  540]='h00000698;  wr_data_rom[  540]='h0000040b;
    rd_cycle[  541] = 1'b0;  wr_cycle[  541] = 1'b1;  addr_rom[  541]='h000002c0;  wr_data_rom[  541]='h00000635;
    rd_cycle[  542] = 1'b0;  wr_cycle[  542] = 1'b1;  addr_rom[  542]='h000003bc;  wr_data_rom[  542]='h000005c0;
    rd_cycle[  543] = 1'b0;  wr_cycle[  543] = 1'b1;  addr_rom[  543]='h00000528;  wr_data_rom[  543]='h000006ae;
    rd_cycle[  544] = 1'b0;  wr_cycle[  544] = 1'b1;  addr_rom[  544]='h00000684;  wr_data_rom[  544]='h000007c3;
    rd_cycle[  545] = 1'b0;  wr_cycle[  545] = 1'b1;  addr_rom[  545]='h000000e0;  wr_data_rom[  545]='h00000633;
    rd_cycle[  546] = 1'b1;  wr_cycle[  546] = 1'b0;  addr_rom[  546]='h00000004;  wr_data_rom[  546]='h00000000;
    rd_cycle[  547] = 1'b0;  wr_cycle[  547] = 1'b1;  addr_rom[  547]='h00000390;  wr_data_rom[  547]='h000007f8;
    rd_cycle[  548] = 1'b0;  wr_cycle[  548] = 1'b1;  addr_rom[  548]='h000004c4;  wr_data_rom[  548]='h00000034;
    rd_cycle[  549] = 1'b0;  wr_cycle[  549] = 1'b1;  addr_rom[  549]='h00000600;  wr_data_rom[  549]='h0000033c;
    rd_cycle[  550] = 1'b1;  wr_cycle[  550] = 1'b0;  addr_rom[  550]='h00000484;  wr_data_rom[  550]='h00000000;
    rd_cycle[  551] = 1'b1;  wr_cycle[  551] = 1'b0;  addr_rom[  551]='h00000210;  wr_data_rom[  551]='h00000000;
    rd_cycle[  552] = 1'b0;  wr_cycle[  552] = 1'b1;  addr_rom[  552]='h000002a4;  wr_data_rom[  552]='h000000d8;
    rd_cycle[  553] = 1'b1;  wr_cycle[  553] = 1'b0;  addr_rom[  553]='h0000060c;  wr_data_rom[  553]='h00000000;
    rd_cycle[  554] = 1'b1;  wr_cycle[  554] = 1'b0;  addr_rom[  554]='h000006e0;  wr_data_rom[  554]='h00000000;
    rd_cycle[  555] = 1'b1;  wr_cycle[  555] = 1'b0;  addr_rom[  555]='h00000044;  wr_data_rom[  555]='h00000000;
    rd_cycle[  556] = 1'b1;  wr_cycle[  556] = 1'b0;  addr_rom[  556]='h00000790;  wr_data_rom[  556]='h00000000;
    rd_cycle[  557] = 1'b1;  wr_cycle[  557] = 1'b0;  addr_rom[  557]='h00000548;  wr_data_rom[  557]='h00000000;
    rd_cycle[  558] = 1'b1;  wr_cycle[  558] = 1'b0;  addr_rom[  558]='h000004b0;  wr_data_rom[  558]='h00000000;
    rd_cycle[  559] = 1'b1;  wr_cycle[  559] = 1'b0;  addr_rom[  559]='h00000498;  wr_data_rom[  559]='h00000000;
    rd_cycle[  560] = 1'b1;  wr_cycle[  560] = 1'b0;  addr_rom[  560]='h0000018c;  wr_data_rom[  560]='h00000000;
    rd_cycle[  561] = 1'b0;  wr_cycle[  561] = 1'b1;  addr_rom[  561]='h000001d8;  wr_data_rom[  561]='h000000f2;
    rd_cycle[  562] = 1'b0;  wr_cycle[  562] = 1'b1;  addr_rom[  562]='h0000073c;  wr_data_rom[  562]='h0000061a;
    rd_cycle[  563] = 1'b0;  wr_cycle[  563] = 1'b1;  addr_rom[  563]='h000004a4;  wr_data_rom[  563]='h000005e7;
    rd_cycle[  564] = 1'b0;  wr_cycle[  564] = 1'b1;  addr_rom[  564]='h000000bc;  wr_data_rom[  564]='h000007c2;
    rd_cycle[  565] = 1'b0;  wr_cycle[  565] = 1'b1;  addr_rom[  565]='h00000098;  wr_data_rom[  565]='h00000432;
    rd_cycle[  566] = 1'b0;  wr_cycle[  566] = 1'b1;  addr_rom[  566]='h00000028;  wr_data_rom[  566]='h00000620;
    rd_cycle[  567] = 1'b1;  wr_cycle[  567] = 1'b0;  addr_rom[  567]='h00000714;  wr_data_rom[  567]='h00000000;
    rd_cycle[  568] = 1'b0;  wr_cycle[  568] = 1'b1;  addr_rom[  568]='h000000a4;  wr_data_rom[  568]='h0000023d;
    rd_cycle[  569] = 1'b0;  wr_cycle[  569] = 1'b1;  addr_rom[  569]='h00000670;  wr_data_rom[  569]='h0000044d;
    rd_cycle[  570] = 1'b1;  wr_cycle[  570] = 1'b0;  addr_rom[  570]='h0000026c;  wr_data_rom[  570]='h00000000;
    rd_cycle[  571] = 1'b0;  wr_cycle[  571] = 1'b1;  addr_rom[  571]='h00000784;  wr_data_rom[  571]='h00000278;
    rd_cycle[  572] = 1'b1;  wr_cycle[  572] = 1'b0;  addr_rom[  572]='h000000d8;  wr_data_rom[  572]='h00000000;
    rd_cycle[  573] = 1'b1;  wr_cycle[  573] = 1'b0;  addr_rom[  573]='h00000368;  wr_data_rom[  573]='h00000000;
    rd_cycle[  574] = 1'b1;  wr_cycle[  574] = 1'b0;  addr_rom[  574]='h000002f4;  wr_data_rom[  574]='h00000000;
    rd_cycle[  575] = 1'b1;  wr_cycle[  575] = 1'b0;  addr_rom[  575]='h00000230;  wr_data_rom[  575]='h00000000;
    rd_cycle[  576] = 1'b1;  wr_cycle[  576] = 1'b0;  addr_rom[  576]='h00000574;  wr_data_rom[  576]='h00000000;
    rd_cycle[  577] = 1'b1;  wr_cycle[  577] = 1'b0;  addr_rom[  577]='h00000208;  wr_data_rom[  577]='h00000000;
    rd_cycle[  578] = 1'b1;  wr_cycle[  578] = 1'b0;  addr_rom[  578]='h00000328;  wr_data_rom[  578]='h00000000;
    rd_cycle[  579] = 1'b0;  wr_cycle[  579] = 1'b1;  addr_rom[  579]='h00000500;  wr_data_rom[  579]='h000007e9;
    rd_cycle[  580] = 1'b0;  wr_cycle[  580] = 1'b1;  addr_rom[  580]='h000001f0;  wr_data_rom[  580]='h000007f0;
    rd_cycle[  581] = 1'b0;  wr_cycle[  581] = 1'b1;  addr_rom[  581]='h00000418;  wr_data_rom[  581]='h000005df;
    rd_cycle[  582] = 1'b0;  wr_cycle[  582] = 1'b1;  addr_rom[  582]='h00000350;  wr_data_rom[  582]='h00000777;
    rd_cycle[  583] = 1'b1;  wr_cycle[  583] = 1'b0;  addr_rom[  583]='h00000088;  wr_data_rom[  583]='h00000000;
    rd_cycle[  584] = 1'b0;  wr_cycle[  584] = 1'b1;  addr_rom[  584]='h0000060c;  wr_data_rom[  584]='h00000266;
    rd_cycle[  585] = 1'b1;  wr_cycle[  585] = 1'b0;  addr_rom[  585]='h0000024c;  wr_data_rom[  585]='h00000000;
    rd_cycle[  586] = 1'b0;  wr_cycle[  586] = 1'b1;  addr_rom[  586]='h00000000;  wr_data_rom[  586]='h00000303;
    rd_cycle[  587] = 1'b0;  wr_cycle[  587] = 1'b1;  addr_rom[  587]='h000002d8;  wr_data_rom[  587]='h0000063f;
    rd_cycle[  588] = 1'b1;  wr_cycle[  588] = 1'b0;  addr_rom[  588]='h000005cc;  wr_data_rom[  588]='h00000000;
    rd_cycle[  589] = 1'b0;  wr_cycle[  589] = 1'b1;  addr_rom[  589]='h00000124;  wr_data_rom[  589]='h00000057;
    rd_cycle[  590] = 1'b0;  wr_cycle[  590] = 1'b1;  addr_rom[  590]='h00000698;  wr_data_rom[  590]='h00000691;
    rd_cycle[  591] = 1'b1;  wr_cycle[  591] = 1'b0;  addr_rom[  591]='h000001a8;  wr_data_rom[  591]='h00000000;
    rd_cycle[  592] = 1'b0;  wr_cycle[  592] = 1'b1;  addr_rom[  592]='h000002f8;  wr_data_rom[  592]='h0000061e;
    rd_cycle[  593] = 1'b0;  wr_cycle[  593] = 1'b1;  addr_rom[  593]='h00000100;  wr_data_rom[  593]='h000000a9;
    rd_cycle[  594] = 1'b0;  wr_cycle[  594] = 1'b1;  addr_rom[  594]='h0000007c;  wr_data_rom[  594]='h000006b5;
    rd_cycle[  595] = 1'b1;  wr_cycle[  595] = 1'b0;  addr_rom[  595]='h00000734;  wr_data_rom[  595]='h00000000;
    rd_cycle[  596] = 1'b0;  wr_cycle[  596] = 1'b1;  addr_rom[  596]='h000004cc;  wr_data_rom[  596]='h000001dc;
    rd_cycle[  597] = 1'b0;  wr_cycle[  597] = 1'b1;  addr_rom[  597]='h000007d4;  wr_data_rom[  597]='h00000639;
    rd_cycle[  598] = 1'b0;  wr_cycle[  598] = 1'b1;  addr_rom[  598]='h000007d0;  wr_data_rom[  598]='h000000ea;
    rd_cycle[  599] = 1'b0;  wr_cycle[  599] = 1'b1;  addr_rom[  599]='h00000420;  wr_data_rom[  599]='h000007f4;
    rd_cycle[  600] = 1'b0;  wr_cycle[  600] = 1'b1;  addr_rom[  600]='h00000598;  wr_data_rom[  600]='h00000016;
    rd_cycle[  601] = 1'b0;  wr_cycle[  601] = 1'b1;  addr_rom[  601]='h000002a4;  wr_data_rom[  601]='h000001c3;
    rd_cycle[  602] = 1'b1;  wr_cycle[  602] = 1'b0;  addr_rom[  602]='h00000608;  wr_data_rom[  602]='h00000000;
    rd_cycle[  603] = 1'b0;  wr_cycle[  603] = 1'b1;  addr_rom[  603]='h0000061c;  wr_data_rom[  603]='h00000137;
    rd_cycle[  604] = 1'b1;  wr_cycle[  604] = 1'b0;  addr_rom[  604]='h00000560;  wr_data_rom[  604]='h00000000;
    rd_cycle[  605] = 1'b0;  wr_cycle[  605] = 1'b1;  addr_rom[  605]='h000001d4;  wr_data_rom[  605]='h000001a9;
    rd_cycle[  606] = 1'b0;  wr_cycle[  606] = 1'b1;  addr_rom[  606]='h00000370;  wr_data_rom[  606]='h000006e8;
    rd_cycle[  607] = 1'b1;  wr_cycle[  607] = 1'b0;  addr_rom[  607]='h00000344;  wr_data_rom[  607]='h00000000;
    rd_cycle[  608] = 1'b0;  wr_cycle[  608] = 1'b1;  addr_rom[  608]='h000003a8;  wr_data_rom[  608]='h00000724;
    rd_cycle[  609] = 1'b1;  wr_cycle[  609] = 1'b0;  addr_rom[  609]='h000002dc;  wr_data_rom[  609]='h00000000;
    rd_cycle[  610] = 1'b0;  wr_cycle[  610] = 1'b1;  addr_rom[  610]='h000007ac;  wr_data_rom[  610]='h00000764;
    rd_cycle[  611] = 1'b0;  wr_cycle[  611] = 1'b1;  addr_rom[  611]='h00000004;  wr_data_rom[  611]='h000003e6;
    rd_cycle[  612] = 1'b1;  wr_cycle[  612] = 1'b0;  addr_rom[  612]='h000003e8;  wr_data_rom[  612]='h00000000;
    rd_cycle[  613] = 1'b1;  wr_cycle[  613] = 1'b0;  addr_rom[  613]='h000007a0;  wr_data_rom[  613]='h00000000;
    rd_cycle[  614] = 1'b1;  wr_cycle[  614] = 1'b0;  addr_rom[  614]='h00000280;  wr_data_rom[  614]='h00000000;
    rd_cycle[  615] = 1'b1;  wr_cycle[  615] = 1'b0;  addr_rom[  615]='h000000b4;  wr_data_rom[  615]='h00000000;
    rd_cycle[  616] = 1'b0;  wr_cycle[  616] = 1'b1;  addr_rom[  616]='h00000278;  wr_data_rom[  616]='h00000255;
    rd_cycle[  617] = 1'b1;  wr_cycle[  617] = 1'b0;  addr_rom[  617]='h00000350;  wr_data_rom[  617]='h00000000;
    rd_cycle[  618] = 1'b0;  wr_cycle[  618] = 1'b1;  addr_rom[  618]='h000000ac;  wr_data_rom[  618]='h000005d0;
    rd_cycle[  619] = 1'b0;  wr_cycle[  619] = 1'b1;  addr_rom[  619]='h0000023c;  wr_data_rom[  619]='h00000226;
    rd_cycle[  620] = 1'b1;  wr_cycle[  620] = 1'b0;  addr_rom[  620]='h00000274;  wr_data_rom[  620]='h00000000;
    rd_cycle[  621] = 1'b0;  wr_cycle[  621] = 1'b1;  addr_rom[  621]='h000004d4;  wr_data_rom[  621]='h000002fc;
    rd_cycle[  622] = 1'b0;  wr_cycle[  622] = 1'b1;  addr_rom[  622]='h000006ac;  wr_data_rom[  622]='h00000463;
    rd_cycle[  623] = 1'b1;  wr_cycle[  623] = 1'b0;  addr_rom[  623]='h00000320;  wr_data_rom[  623]='h00000000;
    rd_cycle[  624] = 1'b0;  wr_cycle[  624] = 1'b1;  addr_rom[  624]='h00000260;  wr_data_rom[  624]='h00000462;
    rd_cycle[  625] = 1'b1;  wr_cycle[  625] = 1'b0;  addr_rom[  625]='h00000690;  wr_data_rom[  625]='h00000000;
    rd_cycle[  626] = 1'b0;  wr_cycle[  626] = 1'b1;  addr_rom[  626]='h000004f0;  wr_data_rom[  626]='h000006a8;
    rd_cycle[  627] = 1'b0;  wr_cycle[  627] = 1'b1;  addr_rom[  627]='h00000144;  wr_data_rom[  627]='h00000459;
    rd_cycle[  628] = 1'b1;  wr_cycle[  628] = 1'b0;  addr_rom[  628]='h0000013c;  wr_data_rom[  628]='h00000000;
    rd_cycle[  629] = 1'b1;  wr_cycle[  629] = 1'b0;  addr_rom[  629]='h000005e4;  wr_data_rom[  629]='h00000000;
    rd_cycle[  630] = 1'b1;  wr_cycle[  630] = 1'b0;  addr_rom[  630]='h00000374;  wr_data_rom[  630]='h00000000;
    rd_cycle[  631] = 1'b0;  wr_cycle[  631] = 1'b1;  addr_rom[  631]='h00000538;  wr_data_rom[  631]='h00000498;
    rd_cycle[  632] = 1'b0;  wr_cycle[  632] = 1'b1;  addr_rom[  632]='h0000004c;  wr_data_rom[  632]='h000000f2;
    rd_cycle[  633] = 1'b1;  wr_cycle[  633] = 1'b0;  addr_rom[  633]='h00000074;  wr_data_rom[  633]='h00000000;
    rd_cycle[  634] = 1'b1;  wr_cycle[  634] = 1'b0;  addr_rom[  634]='h0000006c;  wr_data_rom[  634]='h00000000;
    rd_cycle[  635] = 1'b0;  wr_cycle[  635] = 1'b1;  addr_rom[  635]='h0000046c;  wr_data_rom[  635]='h00000117;
    rd_cycle[  636] = 1'b1;  wr_cycle[  636] = 1'b0;  addr_rom[  636]='h000000d0;  wr_data_rom[  636]='h00000000;
    rd_cycle[  637] = 1'b1;  wr_cycle[  637] = 1'b0;  addr_rom[  637]='h0000006c;  wr_data_rom[  637]='h00000000;
    rd_cycle[  638] = 1'b0;  wr_cycle[  638] = 1'b1;  addr_rom[  638]='h00000440;  wr_data_rom[  638]='h00000718;
    rd_cycle[  639] = 1'b0;  wr_cycle[  639] = 1'b1;  addr_rom[  639]='h00000624;  wr_data_rom[  639]='h00000140;
    rd_cycle[  640] = 1'b1;  wr_cycle[  640] = 1'b0;  addr_rom[  640]='h000002f4;  wr_data_rom[  640]='h00000000;
    rd_cycle[  641] = 1'b0;  wr_cycle[  641] = 1'b1;  addr_rom[  641]='h00000554;  wr_data_rom[  641]='h000005f1;
    rd_cycle[  642] = 1'b0;  wr_cycle[  642] = 1'b1;  addr_rom[  642]='h000006a8;  wr_data_rom[  642]='h00000398;
    rd_cycle[  643] = 1'b1;  wr_cycle[  643] = 1'b0;  addr_rom[  643]='h000002fc;  wr_data_rom[  643]='h00000000;
    rd_cycle[  644] = 1'b0;  wr_cycle[  644] = 1'b1;  addr_rom[  644]='h000006f0;  wr_data_rom[  644]='h00000002;
    rd_cycle[  645] = 1'b0;  wr_cycle[  645] = 1'b1;  addr_rom[  645]='h000002a8;  wr_data_rom[  645]='h00000214;
    rd_cycle[  646] = 1'b1;  wr_cycle[  646] = 1'b0;  addr_rom[  646]='h000005d0;  wr_data_rom[  646]='h00000000;
    rd_cycle[  647] = 1'b0;  wr_cycle[  647] = 1'b1;  addr_rom[  647]='h00000058;  wr_data_rom[  647]='h00000712;
    rd_cycle[  648] = 1'b1;  wr_cycle[  648] = 1'b0;  addr_rom[  648]='h00000744;  wr_data_rom[  648]='h00000000;
    rd_cycle[  649] = 1'b0;  wr_cycle[  649] = 1'b1;  addr_rom[  649]='h000003f4;  wr_data_rom[  649]='h000005ed;
    rd_cycle[  650] = 1'b1;  wr_cycle[  650] = 1'b0;  addr_rom[  650]='h000005ac;  wr_data_rom[  650]='h00000000;
    rd_cycle[  651] = 1'b0;  wr_cycle[  651] = 1'b1;  addr_rom[  651]='h000003e8;  wr_data_rom[  651]='h0000050f;
    rd_cycle[  652] = 1'b1;  wr_cycle[  652] = 1'b0;  addr_rom[  652]='h00000754;  wr_data_rom[  652]='h00000000;
    rd_cycle[  653] = 1'b0;  wr_cycle[  653] = 1'b1;  addr_rom[  653]='h00000390;  wr_data_rom[  653]='h000006e4;
    rd_cycle[  654] = 1'b0;  wr_cycle[  654] = 1'b1;  addr_rom[  654]='h000003a8;  wr_data_rom[  654]='h00000111;
    rd_cycle[  655] = 1'b1;  wr_cycle[  655] = 1'b0;  addr_rom[  655]='h000005a4;  wr_data_rom[  655]='h00000000;
    rd_cycle[  656] = 1'b0;  wr_cycle[  656] = 1'b1;  addr_rom[  656]='h000002f4;  wr_data_rom[  656]='h00000033;
    rd_cycle[  657] = 1'b1;  wr_cycle[  657] = 1'b0;  addr_rom[  657]='h00000454;  wr_data_rom[  657]='h00000000;
    rd_cycle[  658] = 1'b0;  wr_cycle[  658] = 1'b1;  addr_rom[  658]='h0000009c;  wr_data_rom[  658]='h00000068;
    rd_cycle[  659] = 1'b1;  wr_cycle[  659] = 1'b0;  addr_rom[  659]='h00000394;  wr_data_rom[  659]='h00000000;
    rd_cycle[  660] = 1'b0;  wr_cycle[  660] = 1'b1;  addr_rom[  660]='h000001bc;  wr_data_rom[  660]='h00000241;
    rd_cycle[  661] = 1'b0;  wr_cycle[  661] = 1'b1;  addr_rom[  661]='h000000c8;  wr_data_rom[  661]='h0000011f;
    rd_cycle[  662] = 1'b0;  wr_cycle[  662] = 1'b1;  addr_rom[  662]='h00000458;  wr_data_rom[  662]='h00000537;
    rd_cycle[  663] = 1'b1;  wr_cycle[  663] = 1'b0;  addr_rom[  663]='h000002dc;  wr_data_rom[  663]='h00000000;
    rd_cycle[  664] = 1'b1;  wr_cycle[  664] = 1'b0;  addr_rom[  664]='h000003f0;  wr_data_rom[  664]='h00000000;
    rd_cycle[  665] = 1'b0;  wr_cycle[  665] = 1'b1;  addr_rom[  665]='h000003c0;  wr_data_rom[  665]='h000000b2;
    rd_cycle[  666] = 1'b1;  wr_cycle[  666] = 1'b0;  addr_rom[  666]='h00000498;  wr_data_rom[  666]='h00000000;
    rd_cycle[  667] = 1'b1;  wr_cycle[  667] = 1'b0;  addr_rom[  667]='h00000728;  wr_data_rom[  667]='h00000000;
    rd_cycle[  668] = 1'b1;  wr_cycle[  668] = 1'b0;  addr_rom[  668]='h00000560;  wr_data_rom[  668]='h00000000;
    rd_cycle[  669] = 1'b0;  wr_cycle[  669] = 1'b1;  addr_rom[  669]='h000001cc;  wr_data_rom[  669]='h0000042d;
    rd_cycle[  670] = 1'b1;  wr_cycle[  670] = 1'b0;  addr_rom[  670]='h00000284;  wr_data_rom[  670]='h00000000;
    rd_cycle[  671] = 1'b0;  wr_cycle[  671] = 1'b1;  addr_rom[  671]='h000005bc;  wr_data_rom[  671]='h000003c6;
    rd_cycle[  672] = 1'b0;  wr_cycle[  672] = 1'b1;  addr_rom[  672]='h0000032c;  wr_data_rom[  672]='h0000043d;
    rd_cycle[  673] = 1'b1;  wr_cycle[  673] = 1'b0;  addr_rom[  673]='h000004d0;  wr_data_rom[  673]='h00000000;
    rd_cycle[  674] = 1'b0;  wr_cycle[  674] = 1'b1;  addr_rom[  674]='h000006d4;  wr_data_rom[  674]='h00000153;
    rd_cycle[  675] = 1'b0;  wr_cycle[  675] = 1'b1;  addr_rom[  675]='h000000a4;  wr_data_rom[  675]='h00000290;
    rd_cycle[  676] = 1'b0;  wr_cycle[  676] = 1'b1;  addr_rom[  676]='h00000174;  wr_data_rom[  676]='h00000312;
    rd_cycle[  677] = 1'b0;  wr_cycle[  677] = 1'b1;  addr_rom[  677]='h00000288;  wr_data_rom[  677]='h000004b9;
    rd_cycle[  678] = 1'b0;  wr_cycle[  678] = 1'b1;  addr_rom[  678]='h00000598;  wr_data_rom[  678]='h0000055e;
    rd_cycle[  679] = 1'b0;  wr_cycle[  679] = 1'b1;  addr_rom[  679]='h00000560;  wr_data_rom[  679]='h0000058f;
    rd_cycle[  680] = 1'b0;  wr_cycle[  680] = 1'b1;  addr_rom[  680]='h00000754;  wr_data_rom[  680]='h00000690;
    rd_cycle[  681] = 1'b1;  wr_cycle[  681] = 1'b0;  addr_rom[  681]='h00000318;  wr_data_rom[  681]='h00000000;
    rd_cycle[  682] = 1'b0;  wr_cycle[  682] = 1'b1;  addr_rom[  682]='h00000690;  wr_data_rom[  682]='h000007a7;
    rd_cycle[  683] = 1'b1;  wr_cycle[  683] = 1'b0;  addr_rom[  683]='h00000640;  wr_data_rom[  683]='h00000000;
    rd_cycle[  684] = 1'b1;  wr_cycle[  684] = 1'b0;  addr_rom[  684]='h000002a0;  wr_data_rom[  684]='h00000000;
    rd_cycle[  685] = 1'b1;  wr_cycle[  685] = 1'b0;  addr_rom[  685]='h00000690;  wr_data_rom[  685]='h00000000;
    rd_cycle[  686] = 1'b1;  wr_cycle[  686] = 1'b0;  addr_rom[  686]='h000007d4;  wr_data_rom[  686]='h00000000;
    rd_cycle[  687] = 1'b1;  wr_cycle[  687] = 1'b0;  addr_rom[  687]='h000005b4;  wr_data_rom[  687]='h00000000;
    rd_cycle[  688] = 1'b1;  wr_cycle[  688] = 1'b0;  addr_rom[  688]='h000002c4;  wr_data_rom[  688]='h00000000;
    rd_cycle[  689] = 1'b1;  wr_cycle[  689] = 1'b0;  addr_rom[  689]='h0000062c;  wr_data_rom[  689]='h00000000;
    rd_cycle[  690] = 1'b1;  wr_cycle[  690] = 1'b0;  addr_rom[  690]='h000006f4;  wr_data_rom[  690]='h00000000;
    rd_cycle[  691] = 1'b1;  wr_cycle[  691] = 1'b0;  addr_rom[  691]='h000007b8;  wr_data_rom[  691]='h00000000;
    rd_cycle[  692] = 1'b1;  wr_cycle[  692] = 1'b0;  addr_rom[  692]='h00000734;  wr_data_rom[  692]='h00000000;
    rd_cycle[  693] = 1'b0;  wr_cycle[  693] = 1'b1;  addr_rom[  693]='h00000458;  wr_data_rom[  693]='h000000d1;
    rd_cycle[  694] = 1'b1;  wr_cycle[  694] = 1'b0;  addr_rom[  694]='h00000308;  wr_data_rom[  694]='h00000000;
    rd_cycle[  695] = 1'b0;  wr_cycle[  695] = 1'b1;  addr_rom[  695]='h00000294;  wr_data_rom[  695]='h000002be;
    rd_cycle[  696] = 1'b1;  wr_cycle[  696] = 1'b0;  addr_rom[  696]='h000005b0;  wr_data_rom[  696]='h00000000;
    rd_cycle[  697] = 1'b0;  wr_cycle[  697] = 1'b1;  addr_rom[  697]='h0000057c;  wr_data_rom[  697]='h000002ed;
    rd_cycle[  698] = 1'b0;  wr_cycle[  698] = 1'b1;  addr_rom[  698]='h000002a4;  wr_data_rom[  698]='h0000024b;
    rd_cycle[  699] = 1'b0;  wr_cycle[  699] = 1'b1;  addr_rom[  699]='h000003e8;  wr_data_rom[  699]='h0000039e;
    rd_cycle[  700] = 1'b1;  wr_cycle[  700] = 1'b0;  addr_rom[  700]='h00000690;  wr_data_rom[  700]='h00000000;
    rd_cycle[  701] = 1'b0;  wr_cycle[  701] = 1'b1;  addr_rom[  701]='h00000570;  wr_data_rom[  701]='h000001a3;
    rd_cycle[  702] = 1'b1;  wr_cycle[  702] = 1'b0;  addr_rom[  702]='h000000c0;  wr_data_rom[  702]='h00000000;
    rd_cycle[  703] = 1'b0;  wr_cycle[  703] = 1'b1;  addr_rom[  703]='h0000006c;  wr_data_rom[  703]='h0000075a;
    rd_cycle[  704] = 1'b0;  wr_cycle[  704] = 1'b1;  addr_rom[  704]='h00000068;  wr_data_rom[  704]='h00000730;
    rd_cycle[  705] = 1'b0;  wr_cycle[  705] = 1'b1;  addr_rom[  705]='h00000620;  wr_data_rom[  705]='h00000468;
    rd_cycle[  706] = 1'b1;  wr_cycle[  706] = 1'b0;  addr_rom[  706]='h00000088;  wr_data_rom[  706]='h00000000;
    rd_cycle[  707] = 1'b0;  wr_cycle[  707] = 1'b1;  addr_rom[  707]='h00000640;  wr_data_rom[  707]='h00000786;
    rd_cycle[  708] = 1'b1;  wr_cycle[  708] = 1'b0;  addr_rom[  708]='h000004f8;  wr_data_rom[  708]='h00000000;
    rd_cycle[  709] = 1'b1;  wr_cycle[  709] = 1'b0;  addr_rom[  709]='h00000078;  wr_data_rom[  709]='h00000000;
    rd_cycle[  710] = 1'b0;  wr_cycle[  710] = 1'b1;  addr_rom[  710]='h00000424;  wr_data_rom[  710]='h00000057;
    rd_cycle[  711] = 1'b1;  wr_cycle[  711] = 1'b0;  addr_rom[  711]='h000002a4;  wr_data_rom[  711]='h00000000;
    rd_cycle[  712] = 1'b0;  wr_cycle[  712] = 1'b1;  addr_rom[  712]='h000003c0;  wr_data_rom[  712]='h000005f5;
    rd_cycle[  713] = 1'b0;  wr_cycle[  713] = 1'b1;  addr_rom[  713]='h0000035c;  wr_data_rom[  713]='h00000661;
    rd_cycle[  714] = 1'b0;  wr_cycle[  714] = 1'b1;  addr_rom[  714]='h0000025c;  wr_data_rom[  714]='h000002e3;
    rd_cycle[  715] = 1'b1;  wr_cycle[  715] = 1'b0;  addr_rom[  715]='h00000414;  wr_data_rom[  715]='h00000000;
    rd_cycle[  716] = 1'b1;  wr_cycle[  716] = 1'b0;  addr_rom[  716]='h0000039c;  wr_data_rom[  716]='h00000000;
    rd_cycle[  717] = 1'b1;  wr_cycle[  717] = 1'b0;  addr_rom[  717]='h00000730;  wr_data_rom[  717]='h00000000;
    rd_cycle[  718] = 1'b1;  wr_cycle[  718] = 1'b0;  addr_rom[  718]='h00000320;  wr_data_rom[  718]='h00000000;
    rd_cycle[  719] = 1'b1;  wr_cycle[  719] = 1'b0;  addr_rom[  719]='h00000248;  wr_data_rom[  719]='h00000000;
    rd_cycle[  720] = 1'b0;  wr_cycle[  720] = 1'b1;  addr_rom[  720]='h000001e8;  wr_data_rom[  720]='h000002d7;
    rd_cycle[  721] = 1'b1;  wr_cycle[  721] = 1'b0;  addr_rom[  721]='h000004c8;  wr_data_rom[  721]='h00000000;
    rd_cycle[  722] = 1'b1;  wr_cycle[  722] = 1'b0;  addr_rom[  722]='h000005e8;  wr_data_rom[  722]='h00000000;
    rd_cycle[  723] = 1'b0;  wr_cycle[  723] = 1'b1;  addr_rom[  723]='h0000042c;  wr_data_rom[  723]='h000005aa;
    rd_cycle[  724] = 1'b1;  wr_cycle[  724] = 1'b0;  addr_rom[  724]='h000001d4;  wr_data_rom[  724]='h00000000;
    rd_cycle[  725] = 1'b1;  wr_cycle[  725] = 1'b0;  addr_rom[  725]='h00000088;  wr_data_rom[  725]='h00000000;
    rd_cycle[  726] = 1'b1;  wr_cycle[  726] = 1'b0;  addr_rom[  726]='h00000334;  wr_data_rom[  726]='h00000000;
    rd_cycle[  727] = 1'b1;  wr_cycle[  727] = 1'b0;  addr_rom[  727]='h00000564;  wr_data_rom[  727]='h00000000;
    rd_cycle[  728] = 1'b1;  wr_cycle[  728] = 1'b0;  addr_rom[  728]='h000003d4;  wr_data_rom[  728]='h00000000;
    rd_cycle[  729] = 1'b1;  wr_cycle[  729] = 1'b0;  addr_rom[  729]='h0000043c;  wr_data_rom[  729]='h00000000;
    rd_cycle[  730] = 1'b0;  wr_cycle[  730] = 1'b1;  addr_rom[  730]='h000005b0;  wr_data_rom[  730]='h000002e9;
    rd_cycle[  731] = 1'b0;  wr_cycle[  731] = 1'b1;  addr_rom[  731]='h000007ac;  wr_data_rom[  731]='h000005b5;
    rd_cycle[  732] = 1'b0;  wr_cycle[  732] = 1'b1;  addr_rom[  732]='h000005d8;  wr_data_rom[  732]='h0000036b;
    rd_cycle[  733] = 1'b1;  wr_cycle[  733] = 1'b0;  addr_rom[  733]='h0000019c;  wr_data_rom[  733]='h00000000;
    rd_cycle[  734] = 1'b0;  wr_cycle[  734] = 1'b1;  addr_rom[  734]='h00000658;  wr_data_rom[  734]='h0000065b;
    rd_cycle[  735] = 1'b0;  wr_cycle[  735] = 1'b1;  addr_rom[  735]='h0000004c;  wr_data_rom[  735]='h000006bb;
    rd_cycle[  736] = 1'b1;  wr_cycle[  736] = 1'b0;  addr_rom[  736]='h000006d4;  wr_data_rom[  736]='h00000000;
    rd_cycle[  737] = 1'b1;  wr_cycle[  737] = 1'b0;  addr_rom[  737]='h000004cc;  wr_data_rom[  737]='h00000000;
    rd_cycle[  738] = 1'b1;  wr_cycle[  738] = 1'b0;  addr_rom[  738]='h0000012c;  wr_data_rom[  738]='h00000000;
    rd_cycle[  739] = 1'b0;  wr_cycle[  739] = 1'b1;  addr_rom[  739]='h0000052c;  wr_data_rom[  739]='h00000617;
    rd_cycle[  740] = 1'b0;  wr_cycle[  740] = 1'b1;  addr_rom[  740]='h0000078c;  wr_data_rom[  740]='h000005f6;
    rd_cycle[  741] = 1'b1;  wr_cycle[  741] = 1'b0;  addr_rom[  741]='h00000670;  wr_data_rom[  741]='h00000000;
    rd_cycle[  742] = 1'b0;  wr_cycle[  742] = 1'b1;  addr_rom[  742]='h0000004c;  wr_data_rom[  742]='h0000004a;
    rd_cycle[  743] = 1'b0;  wr_cycle[  743] = 1'b1;  addr_rom[  743]='h00000124;  wr_data_rom[  743]='h000003b3;
    rd_cycle[  744] = 1'b0;  wr_cycle[  744] = 1'b1;  addr_rom[  744]='h00000684;  wr_data_rom[  744]='h000001d8;
    rd_cycle[  745] = 1'b0;  wr_cycle[  745] = 1'b1;  addr_rom[  745]='h000002c8;  wr_data_rom[  745]='h000002d6;
    rd_cycle[  746] = 1'b0;  wr_cycle[  746] = 1'b1;  addr_rom[  746]='h000002c0;  wr_data_rom[  746]='h00000399;
    rd_cycle[  747] = 1'b1;  wr_cycle[  747] = 1'b0;  addr_rom[  747]='h0000001c;  wr_data_rom[  747]='h00000000;
    rd_cycle[  748] = 1'b1;  wr_cycle[  748] = 1'b0;  addr_rom[  748]='h000006d4;  wr_data_rom[  748]='h00000000;
    rd_cycle[  749] = 1'b0;  wr_cycle[  749] = 1'b1;  addr_rom[  749]='h000005e8;  wr_data_rom[  749]='h0000008b;
    rd_cycle[  750] = 1'b1;  wr_cycle[  750] = 1'b0;  addr_rom[  750]='h0000061c;  wr_data_rom[  750]='h00000000;
    rd_cycle[  751] = 1'b1;  wr_cycle[  751] = 1'b0;  addr_rom[  751]='h00000334;  wr_data_rom[  751]='h00000000;
    rd_cycle[  752] = 1'b0;  wr_cycle[  752] = 1'b1;  addr_rom[  752]='h000004a0;  wr_data_rom[  752]='h00000367;
    rd_cycle[  753] = 1'b1;  wr_cycle[  753] = 1'b0;  addr_rom[  753]='h000005d8;  wr_data_rom[  753]='h00000000;
    rd_cycle[  754] = 1'b1;  wr_cycle[  754] = 1'b0;  addr_rom[  754]='h000003f4;  wr_data_rom[  754]='h00000000;
    rd_cycle[  755] = 1'b0;  wr_cycle[  755] = 1'b1;  addr_rom[  755]='h00000780;  wr_data_rom[  755]='h000000bd;
    rd_cycle[  756] = 1'b1;  wr_cycle[  756] = 1'b0;  addr_rom[  756]='h000000c4;  wr_data_rom[  756]='h00000000;
    rd_cycle[  757] = 1'b1;  wr_cycle[  757] = 1'b0;  addr_rom[  757]='h00000228;  wr_data_rom[  757]='h00000000;
    rd_cycle[  758] = 1'b1;  wr_cycle[  758] = 1'b0;  addr_rom[  758]='h00000038;  wr_data_rom[  758]='h00000000;
    rd_cycle[  759] = 1'b0;  wr_cycle[  759] = 1'b1;  addr_rom[  759]='h0000060c;  wr_data_rom[  759]='h000004bb;
    rd_cycle[  760] = 1'b1;  wr_cycle[  760] = 1'b0;  addr_rom[  760]='h00000064;  wr_data_rom[  760]='h00000000;
    rd_cycle[  761] = 1'b0;  wr_cycle[  761] = 1'b1;  addr_rom[  761]='h00000360;  wr_data_rom[  761]='h0000015b;
    rd_cycle[  762] = 1'b1;  wr_cycle[  762] = 1'b0;  addr_rom[  762]='h000000a8;  wr_data_rom[  762]='h00000000;
    rd_cycle[  763] = 1'b0;  wr_cycle[  763] = 1'b1;  addr_rom[  763]='h000003e0;  wr_data_rom[  763]='h0000044a;
    rd_cycle[  764] = 1'b1;  wr_cycle[  764] = 1'b0;  addr_rom[  764]='h00000670;  wr_data_rom[  764]='h00000000;
    rd_cycle[  765] = 1'b1;  wr_cycle[  765] = 1'b0;  addr_rom[  765]='h00000478;  wr_data_rom[  765]='h00000000;
    rd_cycle[  766] = 1'b1;  wr_cycle[  766] = 1'b0;  addr_rom[  766]='h000003e0;  wr_data_rom[  766]='h00000000;
    rd_cycle[  767] = 1'b0;  wr_cycle[  767] = 1'b1;  addr_rom[  767]='h000002ec;  wr_data_rom[  767]='h00000203;
    rd_cycle[  768] = 1'b1;  wr_cycle[  768] = 1'b0;  addr_rom[  768]='h00000794;  wr_data_rom[  768]='h00000000;
    rd_cycle[  769] = 1'b0;  wr_cycle[  769] = 1'b1;  addr_rom[  769]='h000004d8;  wr_data_rom[  769]='h00000785;
    rd_cycle[  770] = 1'b1;  wr_cycle[  770] = 1'b0;  addr_rom[  770]='h000000e4;  wr_data_rom[  770]='h00000000;
    rd_cycle[  771] = 1'b1;  wr_cycle[  771] = 1'b0;  addr_rom[  771]='h000005ac;  wr_data_rom[  771]='h00000000;
    rd_cycle[  772] = 1'b1;  wr_cycle[  772] = 1'b0;  addr_rom[  772]='h00000364;  wr_data_rom[  772]='h00000000;
    rd_cycle[  773] = 1'b0;  wr_cycle[  773] = 1'b1;  addr_rom[  773]='h000003b0;  wr_data_rom[  773]='h000007a3;
    rd_cycle[  774] = 1'b0;  wr_cycle[  774] = 1'b1;  addr_rom[  774]='h00000734;  wr_data_rom[  774]='h00000609;
    rd_cycle[  775] = 1'b1;  wr_cycle[  775] = 1'b0;  addr_rom[  775]='h00000664;  wr_data_rom[  775]='h00000000;
    rd_cycle[  776] = 1'b1;  wr_cycle[  776] = 1'b0;  addr_rom[  776]='h000006ec;  wr_data_rom[  776]='h00000000;
    rd_cycle[  777] = 1'b0;  wr_cycle[  777] = 1'b1;  addr_rom[  777]='h000006c4;  wr_data_rom[  777]='h000001fe;
    rd_cycle[  778] = 1'b0;  wr_cycle[  778] = 1'b1;  addr_rom[  778]='h00000344;  wr_data_rom[  778]='h00000530;
    rd_cycle[  779] = 1'b1;  wr_cycle[  779] = 1'b0;  addr_rom[  779]='h00000244;  wr_data_rom[  779]='h00000000;
    rd_cycle[  780] = 1'b1;  wr_cycle[  780] = 1'b0;  addr_rom[  780]='h000000b8;  wr_data_rom[  780]='h00000000;
    rd_cycle[  781] = 1'b1;  wr_cycle[  781] = 1'b0;  addr_rom[  781]='h00000184;  wr_data_rom[  781]='h00000000;
    rd_cycle[  782] = 1'b0;  wr_cycle[  782] = 1'b1;  addr_rom[  782]='h0000048c;  wr_data_rom[  782]='h00000526;
    rd_cycle[  783] = 1'b1;  wr_cycle[  783] = 1'b0;  addr_rom[  783]='h000003e4;  wr_data_rom[  783]='h00000000;
    rd_cycle[  784] = 1'b1;  wr_cycle[  784] = 1'b0;  addr_rom[  784]='h0000016c;  wr_data_rom[  784]='h00000000;
    rd_cycle[  785] = 1'b0;  wr_cycle[  785] = 1'b1;  addr_rom[  785]='h000003fc;  wr_data_rom[  785]='h00000516;
    rd_cycle[  786] = 1'b1;  wr_cycle[  786] = 1'b0;  addr_rom[  786]='h000001a4;  wr_data_rom[  786]='h00000000;
    rd_cycle[  787] = 1'b0;  wr_cycle[  787] = 1'b1;  addr_rom[  787]='h00000614;  wr_data_rom[  787]='h0000015e;
    rd_cycle[  788] = 1'b1;  wr_cycle[  788] = 1'b0;  addr_rom[  788]='h0000039c;  wr_data_rom[  788]='h00000000;
    rd_cycle[  789] = 1'b1;  wr_cycle[  789] = 1'b0;  addr_rom[  789]='h000002d4;  wr_data_rom[  789]='h00000000;
    rd_cycle[  790] = 1'b1;  wr_cycle[  790] = 1'b0;  addr_rom[  790]='h00000258;  wr_data_rom[  790]='h00000000;
    rd_cycle[  791] = 1'b1;  wr_cycle[  791] = 1'b0;  addr_rom[  791]='h00000280;  wr_data_rom[  791]='h00000000;
    rd_cycle[  792] = 1'b0;  wr_cycle[  792] = 1'b1;  addr_rom[  792]='h000003d0;  wr_data_rom[  792]='h00000196;
    rd_cycle[  793] = 1'b1;  wr_cycle[  793] = 1'b0;  addr_rom[  793]='h00000210;  wr_data_rom[  793]='h00000000;
    rd_cycle[  794] = 1'b0;  wr_cycle[  794] = 1'b1;  addr_rom[  794]='h00000328;  wr_data_rom[  794]='h000005cb;
    rd_cycle[  795] = 1'b0;  wr_cycle[  795] = 1'b1;  addr_rom[  795]='h00000390;  wr_data_rom[  795]='h0000070e;
    rd_cycle[  796] = 1'b0;  wr_cycle[  796] = 1'b1;  addr_rom[  796]='h000000d4;  wr_data_rom[  796]='h000003d0;
    rd_cycle[  797] = 1'b0;  wr_cycle[  797] = 1'b1;  addr_rom[  797]='h00000068;  wr_data_rom[  797]='h00000301;
    rd_cycle[  798] = 1'b1;  wr_cycle[  798] = 1'b0;  addr_rom[  798]='h00000350;  wr_data_rom[  798]='h00000000;
    rd_cycle[  799] = 1'b1;  wr_cycle[  799] = 1'b0;  addr_rom[  799]='h000007a4;  wr_data_rom[  799]='h00000000;
    rd_cycle[  800] = 1'b1;  wr_cycle[  800] = 1'b0;  addr_rom[  800]='h0000061c;  wr_data_rom[  800]='h00000000;
    rd_cycle[  801] = 1'b0;  wr_cycle[  801] = 1'b1;  addr_rom[  801]='h0000012c;  wr_data_rom[  801]='h00000177;
    rd_cycle[  802] = 1'b0;  wr_cycle[  802] = 1'b1;  addr_rom[  802]='h0000042c;  wr_data_rom[  802]='h000006dd;
    rd_cycle[  803] = 1'b1;  wr_cycle[  803] = 1'b0;  addr_rom[  803]='h00000438;  wr_data_rom[  803]='h00000000;
    rd_cycle[  804] = 1'b0;  wr_cycle[  804] = 1'b1;  addr_rom[  804]='h000003bc;  wr_data_rom[  804]='h00000793;
    rd_cycle[  805] = 1'b0;  wr_cycle[  805] = 1'b1;  addr_rom[  805]='h00000038;  wr_data_rom[  805]='h0000070a;
    rd_cycle[  806] = 1'b1;  wr_cycle[  806] = 1'b0;  addr_rom[  806]='h000007cc;  wr_data_rom[  806]='h00000000;
    rd_cycle[  807] = 1'b1;  wr_cycle[  807] = 1'b0;  addr_rom[  807]='h0000076c;  wr_data_rom[  807]='h00000000;
    rd_cycle[  808] = 1'b1;  wr_cycle[  808] = 1'b0;  addr_rom[  808]='h000002fc;  wr_data_rom[  808]='h00000000;
    rd_cycle[  809] = 1'b0;  wr_cycle[  809] = 1'b1;  addr_rom[  809]='h0000055c;  wr_data_rom[  809]='h000007f9;
    rd_cycle[  810] = 1'b1;  wr_cycle[  810] = 1'b0;  addr_rom[  810]='h0000053c;  wr_data_rom[  810]='h00000000;
    rd_cycle[  811] = 1'b0;  wr_cycle[  811] = 1'b1;  addr_rom[  811]='h00000510;  wr_data_rom[  811]='h000001a6;
    rd_cycle[  812] = 1'b0;  wr_cycle[  812] = 1'b1;  addr_rom[  812]='h000006f8;  wr_data_rom[  812]='h0000035d;
    rd_cycle[  813] = 1'b1;  wr_cycle[  813] = 1'b0;  addr_rom[  813]='h000005c4;  wr_data_rom[  813]='h00000000;
    rd_cycle[  814] = 1'b0;  wr_cycle[  814] = 1'b1;  addr_rom[  814]='h00000410;  wr_data_rom[  814]='h00000227;
    rd_cycle[  815] = 1'b1;  wr_cycle[  815] = 1'b0;  addr_rom[  815]='h00000158;  wr_data_rom[  815]='h00000000;
    rd_cycle[  816] = 1'b1;  wr_cycle[  816] = 1'b0;  addr_rom[  816]='h000002b0;  wr_data_rom[  816]='h00000000;
    rd_cycle[  817] = 1'b1;  wr_cycle[  817] = 1'b0;  addr_rom[  817]='h000005dc;  wr_data_rom[  817]='h00000000;
    rd_cycle[  818] = 1'b0;  wr_cycle[  818] = 1'b1;  addr_rom[  818]='h00000204;  wr_data_rom[  818]='h00000424;
    rd_cycle[  819] = 1'b1;  wr_cycle[  819] = 1'b0;  addr_rom[  819]='h00000418;  wr_data_rom[  819]='h00000000;
    rd_cycle[  820] = 1'b1;  wr_cycle[  820] = 1'b0;  addr_rom[  820]='h000003e0;  wr_data_rom[  820]='h00000000;
    rd_cycle[  821] = 1'b0;  wr_cycle[  821] = 1'b1;  addr_rom[  821]='h000007e4;  wr_data_rom[  821]='h000005cf;
    rd_cycle[  822] = 1'b0;  wr_cycle[  822] = 1'b1;  addr_rom[  822]='h0000073c;  wr_data_rom[  822]='h0000062a;
    rd_cycle[  823] = 1'b0;  wr_cycle[  823] = 1'b1;  addr_rom[  823]='h000005bc;  wr_data_rom[  823]='h00000277;
    rd_cycle[  824] = 1'b1;  wr_cycle[  824] = 1'b0;  addr_rom[  824]='h00000598;  wr_data_rom[  824]='h00000000;
    rd_cycle[  825] = 1'b1;  wr_cycle[  825] = 1'b0;  addr_rom[  825]='h00000044;  wr_data_rom[  825]='h00000000;
    rd_cycle[  826] = 1'b1;  wr_cycle[  826] = 1'b0;  addr_rom[  826]='h00000160;  wr_data_rom[  826]='h00000000;
    rd_cycle[  827] = 1'b0;  wr_cycle[  827] = 1'b1;  addr_rom[  827]='h00000048;  wr_data_rom[  827]='h00000405;
    rd_cycle[  828] = 1'b1;  wr_cycle[  828] = 1'b0;  addr_rom[  828]='h000006b8;  wr_data_rom[  828]='h00000000;
    rd_cycle[  829] = 1'b0;  wr_cycle[  829] = 1'b1;  addr_rom[  829]='h00000550;  wr_data_rom[  829]='h0000059e;
    rd_cycle[  830] = 1'b0;  wr_cycle[  830] = 1'b1;  addr_rom[  830]='h00000698;  wr_data_rom[  830]='h0000018b;
    rd_cycle[  831] = 1'b1;  wr_cycle[  831] = 1'b0;  addr_rom[  831]='h000002b4;  wr_data_rom[  831]='h00000000;
    rd_cycle[  832] = 1'b0;  wr_cycle[  832] = 1'b1;  addr_rom[  832]='h000004d4;  wr_data_rom[  832]='h000004ab;
    rd_cycle[  833] = 1'b1;  wr_cycle[  833] = 1'b0;  addr_rom[  833]='h00000598;  wr_data_rom[  833]='h00000000;
    rd_cycle[  834] = 1'b1;  wr_cycle[  834] = 1'b0;  addr_rom[  834]='h000005bc;  wr_data_rom[  834]='h00000000;
    rd_cycle[  835] = 1'b1;  wr_cycle[  835] = 1'b0;  addr_rom[  835]='h00000748;  wr_data_rom[  835]='h00000000;
    rd_cycle[  836] = 1'b1;  wr_cycle[  836] = 1'b0;  addr_rom[  836]='h00000728;  wr_data_rom[  836]='h00000000;
    rd_cycle[  837] = 1'b0;  wr_cycle[  837] = 1'b1;  addr_rom[  837]='h00000670;  wr_data_rom[  837]='h00000713;
    rd_cycle[  838] = 1'b1;  wr_cycle[  838] = 1'b0;  addr_rom[  838]='h000003f4;  wr_data_rom[  838]='h00000000;
    rd_cycle[  839] = 1'b0;  wr_cycle[  839] = 1'b1;  addr_rom[  839]='h00000190;  wr_data_rom[  839]='h000000ec;
    rd_cycle[  840] = 1'b0;  wr_cycle[  840] = 1'b1;  addr_rom[  840]='h00000588;  wr_data_rom[  840]='h000006e5;
    rd_cycle[  841] = 1'b1;  wr_cycle[  841] = 1'b0;  addr_rom[  841]='h000005d4;  wr_data_rom[  841]='h00000000;
    rd_cycle[  842] = 1'b0;  wr_cycle[  842] = 1'b1;  addr_rom[  842]='h00000430;  wr_data_rom[  842]='h00000696;
    rd_cycle[  843] = 1'b1;  wr_cycle[  843] = 1'b0;  addr_rom[  843]='h000004ac;  wr_data_rom[  843]='h00000000;
    rd_cycle[  844] = 1'b0;  wr_cycle[  844] = 1'b1;  addr_rom[  844]='h000004fc;  wr_data_rom[  844]='h00000772;
    rd_cycle[  845] = 1'b0;  wr_cycle[  845] = 1'b1;  addr_rom[  845]='h00000324;  wr_data_rom[  845]='h000003f2;
    rd_cycle[  846] = 1'b1;  wr_cycle[  846] = 1'b0;  addr_rom[  846]='h00000424;  wr_data_rom[  846]='h00000000;
    rd_cycle[  847] = 1'b1;  wr_cycle[  847] = 1'b0;  addr_rom[  847]='h0000075c;  wr_data_rom[  847]='h00000000;
    rd_cycle[  848] = 1'b0;  wr_cycle[  848] = 1'b1;  addr_rom[  848]='h000004ac;  wr_data_rom[  848]='h00000184;
    rd_cycle[  849] = 1'b0;  wr_cycle[  849] = 1'b1;  addr_rom[  849]='h00000774;  wr_data_rom[  849]='h00000388;
    rd_cycle[  850] = 1'b1;  wr_cycle[  850] = 1'b0;  addr_rom[  850]='h000004f8;  wr_data_rom[  850]='h00000000;
    rd_cycle[  851] = 1'b1;  wr_cycle[  851] = 1'b0;  addr_rom[  851]='h000002f0;  wr_data_rom[  851]='h00000000;
    rd_cycle[  852] = 1'b1;  wr_cycle[  852] = 1'b0;  addr_rom[  852]='h000002c0;  wr_data_rom[  852]='h00000000;
    rd_cycle[  853] = 1'b0;  wr_cycle[  853] = 1'b1;  addr_rom[  853]='h0000038c;  wr_data_rom[  853]='h000007ca;
    rd_cycle[  854] = 1'b0;  wr_cycle[  854] = 1'b1;  addr_rom[  854]='h000005f4;  wr_data_rom[  854]='h000004c6;
    rd_cycle[  855] = 1'b0;  wr_cycle[  855] = 1'b1;  addr_rom[  855]='h00000210;  wr_data_rom[  855]='h000001af;
    rd_cycle[  856] = 1'b0;  wr_cycle[  856] = 1'b1;  addr_rom[  856]='h000003f8;  wr_data_rom[  856]='h000000db;
    rd_cycle[  857] = 1'b1;  wr_cycle[  857] = 1'b0;  addr_rom[  857]='h00000224;  wr_data_rom[  857]='h00000000;
    rd_cycle[  858] = 1'b0;  wr_cycle[  858] = 1'b1;  addr_rom[  858]='h00000604;  wr_data_rom[  858]='h0000035a;
    rd_cycle[  859] = 1'b1;  wr_cycle[  859] = 1'b0;  addr_rom[  859]='h00000014;  wr_data_rom[  859]='h00000000;
    rd_cycle[  860] = 1'b0;  wr_cycle[  860] = 1'b1;  addr_rom[  860]='h00000658;  wr_data_rom[  860]='h0000015c;
    rd_cycle[  861] = 1'b1;  wr_cycle[  861] = 1'b0;  addr_rom[  861]='h00000548;  wr_data_rom[  861]='h00000000;
    rd_cycle[  862] = 1'b0;  wr_cycle[  862] = 1'b1;  addr_rom[  862]='h000005a8;  wr_data_rom[  862]='h000004ed;
    rd_cycle[  863] = 1'b0;  wr_cycle[  863] = 1'b1;  addr_rom[  863]='h0000051c;  wr_data_rom[  863]='h000006fa;
    rd_cycle[  864] = 1'b1;  wr_cycle[  864] = 1'b0;  addr_rom[  864]='h00000484;  wr_data_rom[  864]='h00000000;
    rd_cycle[  865] = 1'b0;  wr_cycle[  865] = 1'b1;  addr_rom[  865]='h00000784;  wr_data_rom[  865]='h00000796;
    rd_cycle[  866] = 1'b0;  wr_cycle[  866] = 1'b1;  addr_rom[  866]='h000006cc;  wr_data_rom[  866]='h000003af;
    rd_cycle[  867] = 1'b1;  wr_cycle[  867] = 1'b0;  addr_rom[  867]='h000006ac;  wr_data_rom[  867]='h00000000;
    rd_cycle[  868] = 1'b0;  wr_cycle[  868] = 1'b1;  addr_rom[  868]='h000003c0;  wr_data_rom[  868]='h00000369;
    rd_cycle[  869] = 1'b1;  wr_cycle[  869] = 1'b0;  addr_rom[  869]='h000003cc;  wr_data_rom[  869]='h00000000;
    rd_cycle[  870] = 1'b0;  wr_cycle[  870] = 1'b1;  addr_rom[  870]='h00000764;  wr_data_rom[  870]='h0000049b;
    rd_cycle[  871] = 1'b1;  wr_cycle[  871] = 1'b0;  addr_rom[  871]='h00000238;  wr_data_rom[  871]='h00000000;
    rd_cycle[  872] = 1'b0;  wr_cycle[  872] = 1'b1;  addr_rom[  872]='h00000264;  wr_data_rom[  872]='h000005b4;
    rd_cycle[  873] = 1'b1;  wr_cycle[  873] = 1'b0;  addr_rom[  873]='h000001c4;  wr_data_rom[  873]='h00000000;
    rd_cycle[  874] = 1'b0;  wr_cycle[  874] = 1'b1;  addr_rom[  874]='h00000414;  wr_data_rom[  874]='h00000734;
    rd_cycle[  875] = 1'b1;  wr_cycle[  875] = 1'b0;  addr_rom[  875]='h0000022c;  wr_data_rom[  875]='h00000000;
    rd_cycle[  876] = 1'b1;  wr_cycle[  876] = 1'b0;  addr_rom[  876]='h000007bc;  wr_data_rom[  876]='h00000000;
    rd_cycle[  877] = 1'b0;  wr_cycle[  877] = 1'b1;  addr_rom[  877]='h00000518;  wr_data_rom[  877]='h00000370;
    rd_cycle[  878] = 1'b0;  wr_cycle[  878] = 1'b1;  addr_rom[  878]='h000001b8;  wr_data_rom[  878]='h00000336;
    rd_cycle[  879] = 1'b0;  wr_cycle[  879] = 1'b1;  addr_rom[  879]='h000000d0;  wr_data_rom[  879]='h00000579;
    rd_cycle[  880] = 1'b0;  wr_cycle[  880] = 1'b1;  addr_rom[  880]='h00000058;  wr_data_rom[  880]='h00000288;
    rd_cycle[  881] = 1'b0;  wr_cycle[  881] = 1'b1;  addr_rom[  881]='h00000334;  wr_data_rom[  881]='h00000761;
    rd_cycle[  882] = 1'b0;  wr_cycle[  882] = 1'b1;  addr_rom[  882]='h000004b4;  wr_data_rom[  882]='h00000096;
    rd_cycle[  883] = 1'b0;  wr_cycle[  883] = 1'b1;  addr_rom[  883]='h000007ac;  wr_data_rom[  883]='h000000a0;
    rd_cycle[  884] = 1'b1;  wr_cycle[  884] = 1'b0;  addr_rom[  884]='h000000b8;  wr_data_rom[  884]='h00000000;
    rd_cycle[  885] = 1'b0;  wr_cycle[  885] = 1'b1;  addr_rom[  885]='h00000480;  wr_data_rom[  885]='h000003d5;
    rd_cycle[  886] = 1'b1;  wr_cycle[  886] = 1'b0;  addr_rom[  886]='h00000584;  wr_data_rom[  886]='h00000000;
    rd_cycle[  887] = 1'b0;  wr_cycle[  887] = 1'b1;  addr_rom[  887]='h00000648;  wr_data_rom[  887]='h000006c3;
    rd_cycle[  888] = 1'b0;  wr_cycle[  888] = 1'b1;  addr_rom[  888]='h0000026c;  wr_data_rom[  888]='h0000007f;
    rd_cycle[  889] = 1'b0;  wr_cycle[  889] = 1'b1;  addr_rom[  889]='h0000061c;  wr_data_rom[  889]='h0000000a;
    rd_cycle[  890] = 1'b0;  wr_cycle[  890] = 1'b1;  addr_rom[  890]='h000003dc;  wr_data_rom[  890]='h00000572;
    rd_cycle[  891] = 1'b0;  wr_cycle[  891] = 1'b1;  addr_rom[  891]='h000002ac;  wr_data_rom[  891]='h00000059;
    rd_cycle[  892] = 1'b0;  wr_cycle[  892] = 1'b1;  addr_rom[  892]='h000006cc;  wr_data_rom[  892]='h00000431;
    rd_cycle[  893] = 1'b1;  wr_cycle[  893] = 1'b0;  addr_rom[  893]='h00000058;  wr_data_rom[  893]='h00000000;
    rd_cycle[  894] = 1'b1;  wr_cycle[  894] = 1'b0;  addr_rom[  894]='h000007d8;  wr_data_rom[  894]='h00000000;
    rd_cycle[  895] = 1'b1;  wr_cycle[  895] = 1'b0;  addr_rom[  895]='h00000554;  wr_data_rom[  895]='h00000000;
    rd_cycle[  896] = 1'b0;  wr_cycle[  896] = 1'b1;  addr_rom[  896]='h00000704;  wr_data_rom[  896]='h0000038a;
    rd_cycle[  897] = 1'b1;  wr_cycle[  897] = 1'b0;  addr_rom[  897]='h000004c0;  wr_data_rom[  897]='h00000000;
    rd_cycle[  898] = 1'b0;  wr_cycle[  898] = 1'b1;  addr_rom[  898]='h000002ec;  wr_data_rom[  898]='h00000791;
    rd_cycle[  899] = 1'b0;  wr_cycle[  899] = 1'b1;  addr_rom[  899]='h000003c8;  wr_data_rom[  899]='h0000046d;
    rd_cycle[  900] = 1'b0;  wr_cycle[  900] = 1'b1;  addr_rom[  900]='h00000068;  wr_data_rom[  900]='h00000144;
    rd_cycle[  901] = 1'b1;  wr_cycle[  901] = 1'b0;  addr_rom[  901]='h000002d8;  wr_data_rom[  901]='h00000000;
    rd_cycle[  902] = 1'b0;  wr_cycle[  902] = 1'b1;  addr_rom[  902]='h000000e4;  wr_data_rom[  902]='h00000763;
    rd_cycle[  903] = 1'b0;  wr_cycle[  903] = 1'b1;  addr_rom[  903]='h00000390;  wr_data_rom[  903]='h0000014f;
    rd_cycle[  904] = 1'b1;  wr_cycle[  904] = 1'b0;  addr_rom[  904]='h000003c0;  wr_data_rom[  904]='h00000000;
    rd_cycle[  905] = 1'b0;  wr_cycle[  905] = 1'b1;  addr_rom[  905]='h000006c0;  wr_data_rom[  905]='h00000083;
    rd_cycle[  906] = 1'b1;  wr_cycle[  906] = 1'b0;  addr_rom[  906]='h0000072c;  wr_data_rom[  906]='h00000000;
    rd_cycle[  907] = 1'b0;  wr_cycle[  907] = 1'b1;  addr_rom[  907]='h00000604;  wr_data_rom[  907]='h000003c7;
    rd_cycle[  908] = 1'b1;  wr_cycle[  908] = 1'b0;  addr_rom[  908]='h00000434;  wr_data_rom[  908]='h00000000;
    rd_cycle[  909] = 1'b1;  wr_cycle[  909] = 1'b0;  addr_rom[  909]='h000002fc;  wr_data_rom[  909]='h00000000;
    rd_cycle[  910] = 1'b0;  wr_cycle[  910] = 1'b1;  addr_rom[  910]='h00000408;  wr_data_rom[  910]='h00000050;
    rd_cycle[  911] = 1'b1;  wr_cycle[  911] = 1'b0;  addr_rom[  911]='h000002bc;  wr_data_rom[  911]='h00000000;
    rd_cycle[  912] = 1'b1;  wr_cycle[  912] = 1'b0;  addr_rom[  912]='h000004a0;  wr_data_rom[  912]='h00000000;
    rd_cycle[  913] = 1'b1;  wr_cycle[  913] = 1'b0;  addr_rom[  913]='h00000560;  wr_data_rom[  913]='h00000000;
    rd_cycle[  914] = 1'b1;  wr_cycle[  914] = 1'b0;  addr_rom[  914]='h00000790;  wr_data_rom[  914]='h00000000;
    rd_cycle[  915] = 1'b1;  wr_cycle[  915] = 1'b0;  addr_rom[  915]='h0000010c;  wr_data_rom[  915]='h00000000;
    rd_cycle[  916] = 1'b1;  wr_cycle[  916] = 1'b0;  addr_rom[  916]='h00000228;  wr_data_rom[  916]='h00000000;
    rd_cycle[  917] = 1'b0;  wr_cycle[  917] = 1'b1;  addr_rom[  917]='h000006e8;  wr_data_rom[  917]='h000001f5;
    rd_cycle[  918] = 1'b0;  wr_cycle[  918] = 1'b1;  addr_rom[  918]='h00000330;  wr_data_rom[  918]='h000003cb;
    rd_cycle[  919] = 1'b0;  wr_cycle[  919] = 1'b1;  addr_rom[  919]='h00000238;  wr_data_rom[  919]='h00000530;
    rd_cycle[  920] = 1'b1;  wr_cycle[  920] = 1'b0;  addr_rom[  920]='h000002b0;  wr_data_rom[  920]='h00000000;
    rd_cycle[  921] = 1'b0;  wr_cycle[  921] = 1'b1;  addr_rom[  921]='h00000134;  wr_data_rom[  921]='h00000234;
    rd_cycle[  922] = 1'b0;  wr_cycle[  922] = 1'b1;  addr_rom[  922]='h00000628;  wr_data_rom[  922]='h000004ed;
    rd_cycle[  923] = 1'b1;  wr_cycle[  923] = 1'b0;  addr_rom[  923]='h00000710;  wr_data_rom[  923]='h00000000;
    rd_cycle[  924] = 1'b0;  wr_cycle[  924] = 1'b1;  addr_rom[  924]='h00000498;  wr_data_rom[  924]='h00000182;
    rd_cycle[  925] = 1'b1;  wr_cycle[  925] = 1'b0;  addr_rom[  925]='h000002dc;  wr_data_rom[  925]='h00000000;
    rd_cycle[  926] = 1'b0;  wr_cycle[  926] = 1'b1;  addr_rom[  926]='h000000c4;  wr_data_rom[  926]='h000002c8;
    rd_cycle[  927] = 1'b0;  wr_cycle[  927] = 1'b1;  addr_rom[  927]='h00000068;  wr_data_rom[  927]='h000005fd;
    rd_cycle[  928] = 1'b1;  wr_cycle[  928] = 1'b0;  addr_rom[  928]='h000004ac;  wr_data_rom[  928]='h00000000;
    rd_cycle[  929] = 1'b0;  wr_cycle[  929] = 1'b1;  addr_rom[  929]='h00000014;  wr_data_rom[  929]='h0000064a;
    rd_cycle[  930] = 1'b1;  wr_cycle[  930] = 1'b0;  addr_rom[  930]='h00000450;  wr_data_rom[  930]='h00000000;
    rd_cycle[  931] = 1'b1;  wr_cycle[  931] = 1'b0;  addr_rom[  931]='h000007b4;  wr_data_rom[  931]='h00000000;
    rd_cycle[  932] = 1'b1;  wr_cycle[  932] = 1'b0;  addr_rom[  932]='h00000660;  wr_data_rom[  932]='h00000000;
    rd_cycle[  933] = 1'b1;  wr_cycle[  933] = 1'b0;  addr_rom[  933]='h000003e8;  wr_data_rom[  933]='h00000000;
    rd_cycle[  934] = 1'b1;  wr_cycle[  934] = 1'b0;  addr_rom[  934]='h000002b0;  wr_data_rom[  934]='h00000000;
    rd_cycle[  935] = 1'b0;  wr_cycle[  935] = 1'b1;  addr_rom[  935]='h00000248;  wr_data_rom[  935]='h00000700;
    rd_cycle[  936] = 1'b0;  wr_cycle[  936] = 1'b1;  addr_rom[  936]='h00000184;  wr_data_rom[  936]='h00000430;
    rd_cycle[  937] = 1'b0;  wr_cycle[  937] = 1'b1;  addr_rom[  937]='h000005e0;  wr_data_rom[  937]='h00000279;
    rd_cycle[  938] = 1'b0;  wr_cycle[  938] = 1'b1;  addr_rom[  938]='h000000b4;  wr_data_rom[  938]='h000003ea;
    rd_cycle[  939] = 1'b0;  wr_cycle[  939] = 1'b1;  addr_rom[  939]='h000000d0;  wr_data_rom[  939]='h0000061a;
    rd_cycle[  940] = 1'b0;  wr_cycle[  940] = 1'b1;  addr_rom[  940]='h000007bc;  wr_data_rom[  940]='h000004ef;
    rd_cycle[  941] = 1'b0;  wr_cycle[  941] = 1'b1;  addr_rom[  941]='h0000000c;  wr_data_rom[  941]='h000003bb;
    rd_cycle[  942] = 1'b0;  wr_cycle[  942] = 1'b1;  addr_rom[  942]='h00000054;  wr_data_rom[  942]='h000005dd;
    rd_cycle[  943] = 1'b0;  wr_cycle[  943] = 1'b1;  addr_rom[  943]='h000007e4;  wr_data_rom[  943]='h00000666;
    rd_cycle[  944] = 1'b1;  wr_cycle[  944] = 1'b0;  addr_rom[  944]='h00000650;  wr_data_rom[  944]='h00000000;
    rd_cycle[  945] = 1'b0;  wr_cycle[  945] = 1'b1;  addr_rom[  945]='h0000007c;  wr_data_rom[  945]='h00000251;
    rd_cycle[  946] = 1'b1;  wr_cycle[  946] = 1'b0;  addr_rom[  946]='h0000023c;  wr_data_rom[  946]='h00000000;
    rd_cycle[  947] = 1'b1;  wr_cycle[  947] = 1'b0;  addr_rom[  947]='h000003b0;  wr_data_rom[  947]='h00000000;
    rd_cycle[  948] = 1'b1;  wr_cycle[  948] = 1'b0;  addr_rom[  948]='h00000008;  wr_data_rom[  948]='h00000000;
    rd_cycle[  949] = 1'b0;  wr_cycle[  949] = 1'b1;  addr_rom[  949]='h00000518;  wr_data_rom[  949]='h000001d1;
    rd_cycle[  950] = 1'b1;  wr_cycle[  950] = 1'b0;  addr_rom[  950]='h000006d0;  wr_data_rom[  950]='h00000000;
    rd_cycle[  951] = 1'b1;  wr_cycle[  951] = 1'b0;  addr_rom[  951]='h000002ec;  wr_data_rom[  951]='h00000000;
    rd_cycle[  952] = 1'b0;  wr_cycle[  952] = 1'b1;  addr_rom[  952]='h00000150;  wr_data_rom[  952]='h0000025c;
    rd_cycle[  953] = 1'b1;  wr_cycle[  953] = 1'b0;  addr_rom[  953]='h0000060c;  wr_data_rom[  953]='h00000000;
    rd_cycle[  954] = 1'b1;  wr_cycle[  954] = 1'b0;  addr_rom[  954]='h00000248;  wr_data_rom[  954]='h00000000;
    rd_cycle[  955] = 1'b0;  wr_cycle[  955] = 1'b1;  addr_rom[  955]='h000002b0;  wr_data_rom[  955]='h00000241;
    rd_cycle[  956] = 1'b0;  wr_cycle[  956] = 1'b1;  addr_rom[  956]='h000005d4;  wr_data_rom[  956]='h000003fa;
    rd_cycle[  957] = 1'b1;  wr_cycle[  957] = 1'b0;  addr_rom[  957]='h00000634;  wr_data_rom[  957]='h00000000;
    rd_cycle[  958] = 1'b1;  wr_cycle[  958] = 1'b0;  addr_rom[  958]='h00000020;  wr_data_rom[  958]='h00000000;
    rd_cycle[  959] = 1'b0;  wr_cycle[  959] = 1'b1;  addr_rom[  959]='h0000030c;  wr_data_rom[  959]='h00000712;
    rd_cycle[  960] = 1'b0;  wr_cycle[  960] = 1'b1;  addr_rom[  960]='h000007a8;  wr_data_rom[  960]='h00000771;
    rd_cycle[  961] = 1'b0;  wr_cycle[  961] = 1'b1;  addr_rom[  961]='h000003dc;  wr_data_rom[  961]='h00000221;
    rd_cycle[  962] = 1'b0;  wr_cycle[  962] = 1'b1;  addr_rom[  962]='h00000000;  wr_data_rom[  962]='h000004dd;
    rd_cycle[  963] = 1'b0;  wr_cycle[  963] = 1'b1;  addr_rom[  963]='h000007dc;  wr_data_rom[  963]='h00000138;
    rd_cycle[  964] = 1'b1;  wr_cycle[  964] = 1'b0;  addr_rom[  964]='h00000610;  wr_data_rom[  964]='h00000000;
    rd_cycle[  965] = 1'b1;  wr_cycle[  965] = 1'b0;  addr_rom[  965]='h00000530;  wr_data_rom[  965]='h00000000;
    rd_cycle[  966] = 1'b1;  wr_cycle[  966] = 1'b0;  addr_rom[  966]='h000000e4;  wr_data_rom[  966]='h00000000;
    rd_cycle[  967] = 1'b1;  wr_cycle[  967] = 1'b0;  addr_rom[  967]='h00000020;  wr_data_rom[  967]='h00000000;
    rd_cycle[  968] = 1'b1;  wr_cycle[  968] = 1'b0;  addr_rom[  968]='h000002f4;  wr_data_rom[  968]='h00000000;
    rd_cycle[  969] = 1'b1;  wr_cycle[  969] = 1'b0;  addr_rom[  969]='h00000014;  wr_data_rom[  969]='h00000000;
    rd_cycle[  970] = 1'b1;  wr_cycle[  970] = 1'b0;  addr_rom[  970]='h000002a4;  wr_data_rom[  970]='h00000000;
    rd_cycle[  971] = 1'b0;  wr_cycle[  971] = 1'b1;  addr_rom[  971]='h00000078;  wr_data_rom[  971]='h0000037b;
    rd_cycle[  972] = 1'b1;  wr_cycle[  972] = 1'b0;  addr_rom[  972]='h00000314;  wr_data_rom[  972]='h00000000;
    rd_cycle[  973] = 1'b1;  wr_cycle[  973] = 1'b0;  addr_rom[  973]='h0000068c;  wr_data_rom[  973]='h00000000;
    rd_cycle[  974] = 1'b1;  wr_cycle[  974] = 1'b0;  addr_rom[  974]='h00000294;  wr_data_rom[  974]='h00000000;
    rd_cycle[  975] = 1'b1;  wr_cycle[  975] = 1'b0;  addr_rom[  975]='h0000055c;  wr_data_rom[  975]='h00000000;
    rd_cycle[  976] = 1'b1;  wr_cycle[  976] = 1'b0;  addr_rom[  976]='h00000768;  wr_data_rom[  976]='h00000000;
    rd_cycle[  977] = 1'b0;  wr_cycle[  977] = 1'b1;  addr_rom[  977]='h000001c4;  wr_data_rom[  977]='h0000028a;
    rd_cycle[  978] = 1'b1;  wr_cycle[  978] = 1'b0;  addr_rom[  978]='h000000f8;  wr_data_rom[  978]='h00000000;
    rd_cycle[  979] = 1'b0;  wr_cycle[  979] = 1'b1;  addr_rom[  979]='h00000470;  wr_data_rom[  979]='h000002a9;
    rd_cycle[  980] = 1'b0;  wr_cycle[  980] = 1'b1;  addr_rom[  980]='h000002d0;  wr_data_rom[  980]='h0000005c;
    rd_cycle[  981] = 1'b1;  wr_cycle[  981] = 1'b0;  addr_rom[  981]='h00000244;  wr_data_rom[  981]='h00000000;
    rd_cycle[  982] = 1'b1;  wr_cycle[  982] = 1'b0;  addr_rom[  982]='h000003c8;  wr_data_rom[  982]='h00000000;
    rd_cycle[  983] = 1'b0;  wr_cycle[  983] = 1'b1;  addr_rom[  983]='h00000384;  wr_data_rom[  983]='h000004c0;
    rd_cycle[  984] = 1'b0;  wr_cycle[  984] = 1'b1;  addr_rom[  984]='h00000628;  wr_data_rom[  984]='h0000015f;
    rd_cycle[  985] = 1'b1;  wr_cycle[  985] = 1'b0;  addr_rom[  985]='h00000164;  wr_data_rom[  985]='h00000000;
    rd_cycle[  986] = 1'b0;  wr_cycle[  986] = 1'b1;  addr_rom[  986]='h00000618;  wr_data_rom[  986]='h00000391;
    rd_cycle[  987] = 1'b1;  wr_cycle[  987] = 1'b0;  addr_rom[  987]='h00000038;  wr_data_rom[  987]='h00000000;
    rd_cycle[  988] = 1'b1;  wr_cycle[  988] = 1'b0;  addr_rom[  988]='h00000044;  wr_data_rom[  988]='h00000000;
    rd_cycle[  989] = 1'b0;  wr_cycle[  989] = 1'b1;  addr_rom[  989]='h00000248;  wr_data_rom[  989]='h000000aa;
    rd_cycle[  990] = 1'b1;  wr_cycle[  990] = 1'b0;  addr_rom[  990]='h00000068;  wr_data_rom[  990]='h00000000;
    rd_cycle[  991] = 1'b1;  wr_cycle[  991] = 1'b0;  addr_rom[  991]='h00000314;  wr_data_rom[  991]='h00000000;
    rd_cycle[  992] = 1'b1;  wr_cycle[  992] = 1'b0;  addr_rom[  992]='h000006e4;  wr_data_rom[  992]='h00000000;
    rd_cycle[  993] = 1'b0;  wr_cycle[  993] = 1'b1;  addr_rom[  993]='h000001e4;  wr_data_rom[  993]='h0000004d;
    rd_cycle[  994] = 1'b0;  wr_cycle[  994] = 1'b1;  addr_rom[  994]='h000007d4;  wr_data_rom[  994]='h000006ea;
    rd_cycle[  995] = 1'b0;  wr_cycle[  995] = 1'b1;  addr_rom[  995]='h00000084;  wr_data_rom[  995]='h000003a5;
    rd_cycle[  996] = 1'b1;  wr_cycle[  996] = 1'b0;  addr_rom[  996]='h0000037c;  wr_data_rom[  996]='h00000000;
    rd_cycle[  997] = 1'b0;  wr_cycle[  997] = 1'b1;  addr_rom[  997]='h000007c0;  wr_data_rom[  997]='h0000006c;
    rd_cycle[  998] = 1'b1;  wr_cycle[  998] = 1'b0;  addr_rom[  998]='h000006d4;  wr_data_rom[  998]='h00000000;
    rd_cycle[  999] = 1'b1;  wr_cycle[  999] = 1'b0;  addr_rom[  999]='h00000250;  wr_data_rom[  999]='h00000000;
    rd_cycle[ 1000] = 1'b0;  wr_cycle[ 1000] = 1'b1;  addr_rom[ 1000]='h000002fc;  wr_data_rom[ 1000]='h00000263;
    rd_cycle[ 1001] = 1'b0;  wr_cycle[ 1001] = 1'b1;  addr_rom[ 1001]='h000007ec;  wr_data_rom[ 1001]='h00000628;
    rd_cycle[ 1002] = 1'b1;  wr_cycle[ 1002] = 1'b0;  addr_rom[ 1002]='h00000640;  wr_data_rom[ 1002]='h00000000;
    rd_cycle[ 1003] = 1'b0;  wr_cycle[ 1003] = 1'b1;  addr_rom[ 1003]='h00000448;  wr_data_rom[ 1003]='h0000018e;
    rd_cycle[ 1004] = 1'b0;  wr_cycle[ 1004] = 1'b1;  addr_rom[ 1004]='h00000560;  wr_data_rom[ 1004]='h0000049f;
    rd_cycle[ 1005] = 1'b1;  wr_cycle[ 1005] = 1'b0;  addr_rom[ 1005]='h000002d0;  wr_data_rom[ 1005]='h00000000;
    rd_cycle[ 1006] = 1'b1;  wr_cycle[ 1006] = 1'b0;  addr_rom[ 1006]='h00000664;  wr_data_rom[ 1006]='h00000000;
    rd_cycle[ 1007] = 1'b1;  wr_cycle[ 1007] = 1'b0;  addr_rom[ 1007]='h0000015c;  wr_data_rom[ 1007]='h00000000;
    rd_cycle[ 1008] = 1'b0;  wr_cycle[ 1008] = 1'b1;  addr_rom[ 1008]='h00000400;  wr_data_rom[ 1008]='h00000078;
    rd_cycle[ 1009] = 1'b1;  wr_cycle[ 1009] = 1'b0;  addr_rom[ 1009]='h00000598;  wr_data_rom[ 1009]='h00000000;
    rd_cycle[ 1010] = 1'b1;  wr_cycle[ 1010] = 1'b0;  addr_rom[ 1010]='h00000620;  wr_data_rom[ 1010]='h00000000;
    rd_cycle[ 1011] = 1'b1;  wr_cycle[ 1011] = 1'b0;  addr_rom[ 1011]='h00000470;  wr_data_rom[ 1011]='h00000000;
    rd_cycle[ 1012] = 1'b0;  wr_cycle[ 1012] = 1'b1;  addr_rom[ 1012]='h00000698;  wr_data_rom[ 1012]='h00000683;
    rd_cycle[ 1013] = 1'b0;  wr_cycle[ 1013] = 1'b1;  addr_rom[ 1013]='h00000498;  wr_data_rom[ 1013]='h00000431;
    rd_cycle[ 1014] = 1'b1;  wr_cycle[ 1014] = 1'b0;  addr_rom[ 1014]='h0000024c;  wr_data_rom[ 1014]='h00000000;
    rd_cycle[ 1015] = 1'b0;  wr_cycle[ 1015] = 1'b1;  addr_rom[ 1015]='h000003b8;  wr_data_rom[ 1015]='h00000142;
    rd_cycle[ 1016] = 1'b0;  wr_cycle[ 1016] = 1'b1;  addr_rom[ 1016]='h00000484;  wr_data_rom[ 1016]='h00000193;
    rd_cycle[ 1017] = 1'b1;  wr_cycle[ 1017] = 1'b0;  addr_rom[ 1017]='h000006b0;  wr_data_rom[ 1017]='h00000000;
    rd_cycle[ 1018] = 1'b0;  wr_cycle[ 1018] = 1'b1;  addr_rom[ 1018]='h000005f0;  wr_data_rom[ 1018]='h000006c8;
    rd_cycle[ 1019] = 1'b1;  wr_cycle[ 1019] = 1'b0;  addr_rom[ 1019]='h00000260;  wr_data_rom[ 1019]='h00000000;
    rd_cycle[ 1020] = 1'b0;  wr_cycle[ 1020] = 1'b1;  addr_rom[ 1020]='h00000694;  wr_data_rom[ 1020]='h00000521;
    rd_cycle[ 1021] = 1'b1;  wr_cycle[ 1021] = 1'b0;  addr_rom[ 1021]='h000007a0;  wr_data_rom[ 1021]='h00000000;
    rd_cycle[ 1022] = 1'b1;  wr_cycle[ 1022] = 1'b0;  addr_rom[ 1022]='h00000188;  wr_data_rom[ 1022]='h00000000;
    rd_cycle[ 1023] = 1'b1;  wr_cycle[ 1023] = 1'b0;  addr_rom[ 1023]='h000006a0;  wr_data_rom[ 1023]='h00000000;
    rd_cycle[ 1024] = 1'b1;  wr_cycle[ 1024] = 1'b0;  addr_rom[ 1024]='h0000048c;  wr_data_rom[ 1024]='h00000000;
    rd_cycle[ 1025] = 1'b0;  wr_cycle[ 1025] = 1'b1;  addr_rom[ 1025]='h000004a0;  wr_data_rom[ 1025]='h00000458;
    rd_cycle[ 1026] = 1'b0;  wr_cycle[ 1026] = 1'b1;  addr_rom[ 1026]='h0000006c;  wr_data_rom[ 1026]='h000006ae;
    rd_cycle[ 1027] = 1'b0;  wr_cycle[ 1027] = 1'b1;  addr_rom[ 1027]='h000003a4;  wr_data_rom[ 1027]='h0000017a;
    rd_cycle[ 1028] = 1'b0;  wr_cycle[ 1028] = 1'b1;  addr_rom[ 1028]='h0000019c;  wr_data_rom[ 1028]='h000000da;
    rd_cycle[ 1029] = 1'b0;  wr_cycle[ 1029] = 1'b1;  addr_rom[ 1029]='h00000070;  wr_data_rom[ 1029]='h0000049a;
    rd_cycle[ 1030] = 1'b0;  wr_cycle[ 1030] = 1'b1;  addr_rom[ 1030]='h000000f8;  wr_data_rom[ 1030]='h000004a0;
    rd_cycle[ 1031] = 1'b1;  wr_cycle[ 1031] = 1'b0;  addr_rom[ 1031]='h000006dc;  wr_data_rom[ 1031]='h00000000;
    rd_cycle[ 1032] = 1'b0;  wr_cycle[ 1032] = 1'b1;  addr_rom[ 1032]='h00000768;  wr_data_rom[ 1032]='h00000640;
    rd_cycle[ 1033] = 1'b0;  wr_cycle[ 1033] = 1'b1;  addr_rom[ 1033]='h00000038;  wr_data_rom[ 1033]='h000001a3;
    rd_cycle[ 1034] = 1'b0;  wr_cycle[ 1034] = 1'b1;  addr_rom[ 1034]='h000006f4;  wr_data_rom[ 1034]='h000005e8;
    rd_cycle[ 1035] = 1'b0;  wr_cycle[ 1035] = 1'b1;  addr_rom[ 1035]='h00000588;  wr_data_rom[ 1035]='h000006b7;
    rd_cycle[ 1036] = 1'b0;  wr_cycle[ 1036] = 1'b1;  addr_rom[ 1036]='h000004ec;  wr_data_rom[ 1036]='h000001e2;
    rd_cycle[ 1037] = 1'b1;  wr_cycle[ 1037] = 1'b0;  addr_rom[ 1037]='h00000410;  wr_data_rom[ 1037]='h00000000;
    rd_cycle[ 1038] = 1'b1;  wr_cycle[ 1038] = 1'b0;  addr_rom[ 1038]='h000002a0;  wr_data_rom[ 1038]='h00000000;
    rd_cycle[ 1039] = 1'b0;  wr_cycle[ 1039] = 1'b1;  addr_rom[ 1039]='h000005ec;  wr_data_rom[ 1039]='h00000486;
    rd_cycle[ 1040] = 1'b0;  wr_cycle[ 1040] = 1'b1;  addr_rom[ 1040]='h000003ec;  wr_data_rom[ 1040]='h00000210;
    rd_cycle[ 1041] = 1'b1;  wr_cycle[ 1041] = 1'b0;  addr_rom[ 1041]='h00000748;  wr_data_rom[ 1041]='h00000000;
    rd_cycle[ 1042] = 1'b1;  wr_cycle[ 1042] = 1'b0;  addr_rom[ 1042]='h0000061c;  wr_data_rom[ 1042]='h00000000;
    rd_cycle[ 1043] = 1'b1;  wr_cycle[ 1043] = 1'b0;  addr_rom[ 1043]='h000000f8;  wr_data_rom[ 1043]='h00000000;
    rd_cycle[ 1044] = 1'b0;  wr_cycle[ 1044] = 1'b1;  addr_rom[ 1044]='h0000061c;  wr_data_rom[ 1044]='h00000413;
    rd_cycle[ 1045] = 1'b0;  wr_cycle[ 1045] = 1'b1;  addr_rom[ 1045]='h0000021c;  wr_data_rom[ 1045]='h00000635;
    rd_cycle[ 1046] = 1'b0;  wr_cycle[ 1046] = 1'b1;  addr_rom[ 1046]='h00000078;  wr_data_rom[ 1046]='h000006ca;
    rd_cycle[ 1047] = 1'b1;  wr_cycle[ 1047] = 1'b0;  addr_rom[ 1047]='h000005a4;  wr_data_rom[ 1047]='h00000000;
    rd_cycle[ 1048] = 1'b0;  wr_cycle[ 1048] = 1'b1;  addr_rom[ 1048]='h000005c0;  wr_data_rom[ 1048]='h00000581;
    rd_cycle[ 1049] = 1'b1;  wr_cycle[ 1049] = 1'b0;  addr_rom[ 1049]='h00000364;  wr_data_rom[ 1049]='h00000000;
    rd_cycle[ 1050] = 1'b0;  wr_cycle[ 1050] = 1'b1;  addr_rom[ 1050]='h00000168;  wr_data_rom[ 1050]='h000000f3;
    rd_cycle[ 1051] = 1'b0;  wr_cycle[ 1051] = 1'b1;  addr_rom[ 1051]='h00000674;  wr_data_rom[ 1051]='h00000761;
    rd_cycle[ 1052] = 1'b0;  wr_cycle[ 1052] = 1'b1;  addr_rom[ 1052]='h00000570;  wr_data_rom[ 1052]='h000006c7;
    rd_cycle[ 1053] = 1'b0;  wr_cycle[ 1053] = 1'b1;  addr_rom[ 1053]='h000006dc;  wr_data_rom[ 1053]='h000000c1;
    rd_cycle[ 1054] = 1'b0;  wr_cycle[ 1054] = 1'b1;  addr_rom[ 1054]='h000007a8;  wr_data_rom[ 1054]='h000003e1;
    rd_cycle[ 1055] = 1'b0;  wr_cycle[ 1055] = 1'b1;  addr_rom[ 1055]='h00000118;  wr_data_rom[ 1055]='h000004a9;
    rd_cycle[ 1056] = 1'b1;  wr_cycle[ 1056] = 1'b0;  addr_rom[ 1056]='h000005d4;  wr_data_rom[ 1056]='h00000000;
    rd_cycle[ 1057] = 1'b0;  wr_cycle[ 1057] = 1'b1;  addr_rom[ 1057]='h000005d4;  wr_data_rom[ 1057]='h00000269;
    rd_cycle[ 1058] = 1'b0;  wr_cycle[ 1058] = 1'b1;  addr_rom[ 1058]='h000006d0;  wr_data_rom[ 1058]='h000006da;
    rd_cycle[ 1059] = 1'b1;  wr_cycle[ 1059] = 1'b0;  addr_rom[ 1059]='h00000714;  wr_data_rom[ 1059]='h00000000;
    rd_cycle[ 1060] = 1'b0;  wr_cycle[ 1060] = 1'b1;  addr_rom[ 1060]='h000005cc;  wr_data_rom[ 1060]='h00000472;
    rd_cycle[ 1061] = 1'b1;  wr_cycle[ 1061] = 1'b0;  addr_rom[ 1061]='h00000678;  wr_data_rom[ 1061]='h00000000;
    rd_cycle[ 1062] = 1'b0;  wr_cycle[ 1062] = 1'b1;  addr_rom[ 1062]='h000007e0;  wr_data_rom[ 1062]='h0000052f;
    rd_cycle[ 1063] = 1'b0;  wr_cycle[ 1063] = 1'b1;  addr_rom[ 1063]='h000001f4;  wr_data_rom[ 1063]='h0000010b;
    rd_cycle[ 1064] = 1'b0;  wr_cycle[ 1064] = 1'b1;  addr_rom[ 1064]='h00000534;  wr_data_rom[ 1064]='h00000727;
    rd_cycle[ 1065] = 1'b0;  wr_cycle[ 1065] = 1'b1;  addr_rom[ 1065]='h00000230;  wr_data_rom[ 1065]='h000007a8;
    rd_cycle[ 1066] = 1'b1;  wr_cycle[ 1066] = 1'b0;  addr_rom[ 1066]='h000007d4;  wr_data_rom[ 1066]='h00000000;
    rd_cycle[ 1067] = 1'b1;  wr_cycle[ 1067] = 1'b0;  addr_rom[ 1067]='h000003f4;  wr_data_rom[ 1067]='h00000000;
    rd_cycle[ 1068] = 1'b1;  wr_cycle[ 1068] = 1'b0;  addr_rom[ 1068]='h00000244;  wr_data_rom[ 1068]='h00000000;
    rd_cycle[ 1069] = 1'b1;  wr_cycle[ 1069] = 1'b0;  addr_rom[ 1069]='h000000fc;  wr_data_rom[ 1069]='h00000000;
    rd_cycle[ 1070] = 1'b1;  wr_cycle[ 1070] = 1'b0;  addr_rom[ 1070]='h00000788;  wr_data_rom[ 1070]='h00000000;
    rd_cycle[ 1071] = 1'b1;  wr_cycle[ 1071] = 1'b0;  addr_rom[ 1071]='h000006c4;  wr_data_rom[ 1071]='h00000000;
    rd_cycle[ 1072] = 1'b1;  wr_cycle[ 1072] = 1'b0;  addr_rom[ 1072]='h000006fc;  wr_data_rom[ 1072]='h00000000;
    rd_cycle[ 1073] = 1'b0;  wr_cycle[ 1073] = 1'b1;  addr_rom[ 1073]='h0000062c;  wr_data_rom[ 1073]='h0000043b;
    rd_cycle[ 1074] = 1'b0;  wr_cycle[ 1074] = 1'b1;  addr_rom[ 1074]='h00000160;  wr_data_rom[ 1074]='h00000519;
    rd_cycle[ 1075] = 1'b0;  wr_cycle[ 1075] = 1'b1;  addr_rom[ 1075]='h000001ec;  wr_data_rom[ 1075]='h00000781;
    rd_cycle[ 1076] = 1'b1;  wr_cycle[ 1076] = 1'b0;  addr_rom[ 1076]='h000003bc;  wr_data_rom[ 1076]='h00000000;
    rd_cycle[ 1077] = 1'b1;  wr_cycle[ 1077] = 1'b0;  addr_rom[ 1077]='h000001dc;  wr_data_rom[ 1077]='h00000000;
    rd_cycle[ 1078] = 1'b1;  wr_cycle[ 1078] = 1'b0;  addr_rom[ 1078]='h00000764;  wr_data_rom[ 1078]='h00000000;
    rd_cycle[ 1079] = 1'b0;  wr_cycle[ 1079] = 1'b1;  addr_rom[ 1079]='h0000057c;  wr_data_rom[ 1079]='h00000176;
    rd_cycle[ 1080] = 1'b0;  wr_cycle[ 1080] = 1'b1;  addr_rom[ 1080]='h00000380;  wr_data_rom[ 1080]='h0000023a;
    rd_cycle[ 1081] = 1'b0;  wr_cycle[ 1081] = 1'b1;  addr_rom[ 1081]='h0000064c;  wr_data_rom[ 1081]='h0000021f;
    rd_cycle[ 1082] = 1'b1;  wr_cycle[ 1082] = 1'b0;  addr_rom[ 1082]='h000000e0;  wr_data_rom[ 1082]='h00000000;
    rd_cycle[ 1083] = 1'b1;  wr_cycle[ 1083] = 1'b0;  addr_rom[ 1083]='h00000238;  wr_data_rom[ 1083]='h00000000;
    rd_cycle[ 1084] = 1'b0;  wr_cycle[ 1084] = 1'b1;  addr_rom[ 1084]='h000002f4;  wr_data_rom[ 1084]='h0000038c;
    rd_cycle[ 1085] = 1'b1;  wr_cycle[ 1085] = 1'b0;  addr_rom[ 1085]='h00000124;  wr_data_rom[ 1085]='h00000000;
    rd_cycle[ 1086] = 1'b1;  wr_cycle[ 1086] = 1'b0;  addr_rom[ 1086]='h00000734;  wr_data_rom[ 1086]='h00000000;
    rd_cycle[ 1087] = 1'b1;  wr_cycle[ 1087] = 1'b0;  addr_rom[ 1087]='h000002bc;  wr_data_rom[ 1087]='h00000000;
    rd_cycle[ 1088] = 1'b1;  wr_cycle[ 1088] = 1'b0;  addr_rom[ 1088]='h000002c4;  wr_data_rom[ 1088]='h00000000;
    rd_cycle[ 1089] = 1'b0;  wr_cycle[ 1089] = 1'b1;  addr_rom[ 1089]='h000006bc;  wr_data_rom[ 1089]='h0000043d;
    rd_cycle[ 1090] = 1'b1;  wr_cycle[ 1090] = 1'b0;  addr_rom[ 1090]='h000002d4;  wr_data_rom[ 1090]='h00000000;
    rd_cycle[ 1091] = 1'b1;  wr_cycle[ 1091] = 1'b0;  addr_rom[ 1091]='h00000708;  wr_data_rom[ 1091]='h00000000;
    rd_cycle[ 1092] = 1'b0;  wr_cycle[ 1092] = 1'b1;  addr_rom[ 1092]='h0000010c;  wr_data_rom[ 1092]='h0000027c;
    rd_cycle[ 1093] = 1'b0;  wr_cycle[ 1093] = 1'b1;  addr_rom[ 1093]='h00000698;  wr_data_rom[ 1093]='h00000617;
    rd_cycle[ 1094] = 1'b0;  wr_cycle[ 1094] = 1'b1;  addr_rom[ 1094]='h00000050;  wr_data_rom[ 1094]='h000002f7;
    rd_cycle[ 1095] = 1'b0;  wr_cycle[ 1095] = 1'b1;  addr_rom[ 1095]='h00000670;  wr_data_rom[ 1095]='h000002ce;
    rd_cycle[ 1096] = 1'b0;  wr_cycle[ 1096] = 1'b1;  addr_rom[ 1096]='h000006b0;  wr_data_rom[ 1096]='h00000240;
    rd_cycle[ 1097] = 1'b0;  wr_cycle[ 1097] = 1'b1;  addr_rom[ 1097]='h000002f4;  wr_data_rom[ 1097]='h000003c5;
    rd_cycle[ 1098] = 1'b1;  wr_cycle[ 1098] = 1'b0;  addr_rom[ 1098]='h00000780;  wr_data_rom[ 1098]='h00000000;
    rd_cycle[ 1099] = 1'b0;  wr_cycle[ 1099] = 1'b1;  addr_rom[ 1099]='h00000204;  wr_data_rom[ 1099]='h00000414;
    rd_cycle[ 1100] = 1'b1;  wr_cycle[ 1100] = 1'b0;  addr_rom[ 1100]='h000005bc;  wr_data_rom[ 1100]='h00000000;
    rd_cycle[ 1101] = 1'b0;  wr_cycle[ 1101] = 1'b1;  addr_rom[ 1101]='h000006f8;  wr_data_rom[ 1101]='h000007a2;
    rd_cycle[ 1102] = 1'b1;  wr_cycle[ 1102] = 1'b0;  addr_rom[ 1102]='h000001dc;  wr_data_rom[ 1102]='h00000000;
    rd_cycle[ 1103] = 1'b0;  wr_cycle[ 1103] = 1'b1;  addr_rom[ 1103]='h000006fc;  wr_data_rom[ 1103]='h00000123;
    rd_cycle[ 1104] = 1'b1;  wr_cycle[ 1104] = 1'b0;  addr_rom[ 1104]='h00000460;  wr_data_rom[ 1104]='h00000000;
    rd_cycle[ 1105] = 1'b1;  wr_cycle[ 1105] = 1'b0;  addr_rom[ 1105]='h000001c4;  wr_data_rom[ 1105]='h00000000;
    rd_cycle[ 1106] = 1'b1;  wr_cycle[ 1106] = 1'b0;  addr_rom[ 1106]='h00000038;  wr_data_rom[ 1106]='h00000000;
    rd_cycle[ 1107] = 1'b1;  wr_cycle[ 1107] = 1'b0;  addr_rom[ 1107]='h00000078;  wr_data_rom[ 1107]='h00000000;
    rd_cycle[ 1108] = 1'b1;  wr_cycle[ 1108] = 1'b0;  addr_rom[ 1108]='h00000578;  wr_data_rom[ 1108]='h00000000;
    rd_cycle[ 1109] = 1'b1;  wr_cycle[ 1109] = 1'b0;  addr_rom[ 1109]='h00000448;  wr_data_rom[ 1109]='h00000000;
    rd_cycle[ 1110] = 1'b0;  wr_cycle[ 1110] = 1'b1;  addr_rom[ 1110]='h00000328;  wr_data_rom[ 1110]='h000000de;
    rd_cycle[ 1111] = 1'b0;  wr_cycle[ 1111] = 1'b1;  addr_rom[ 1111]='h00000048;  wr_data_rom[ 1111]='h000000b2;
    rd_cycle[ 1112] = 1'b1;  wr_cycle[ 1112] = 1'b0;  addr_rom[ 1112]='h000000a4;  wr_data_rom[ 1112]='h00000000;
    rd_cycle[ 1113] = 1'b0;  wr_cycle[ 1113] = 1'b1;  addr_rom[ 1113]='h00000104;  wr_data_rom[ 1113]='h0000069a;
    rd_cycle[ 1114] = 1'b0;  wr_cycle[ 1114] = 1'b1;  addr_rom[ 1114]='h00000614;  wr_data_rom[ 1114]='h00000115;
    rd_cycle[ 1115] = 1'b0;  wr_cycle[ 1115] = 1'b1;  addr_rom[ 1115]='h00000504;  wr_data_rom[ 1115]='h000000b8;
    rd_cycle[ 1116] = 1'b1;  wr_cycle[ 1116] = 1'b0;  addr_rom[ 1116]='h000000a0;  wr_data_rom[ 1116]='h00000000;
    rd_cycle[ 1117] = 1'b0;  wr_cycle[ 1117] = 1'b1;  addr_rom[ 1117]='h000007bc;  wr_data_rom[ 1117]='h00000595;
    rd_cycle[ 1118] = 1'b1;  wr_cycle[ 1118] = 1'b0;  addr_rom[ 1118]='h0000040c;  wr_data_rom[ 1118]='h00000000;
    rd_cycle[ 1119] = 1'b1;  wr_cycle[ 1119] = 1'b0;  addr_rom[ 1119]='h00000158;  wr_data_rom[ 1119]='h00000000;
    rd_cycle[ 1120] = 1'b1;  wr_cycle[ 1120] = 1'b0;  addr_rom[ 1120]='h000006c0;  wr_data_rom[ 1120]='h00000000;
    rd_cycle[ 1121] = 1'b1;  wr_cycle[ 1121] = 1'b0;  addr_rom[ 1121]='h00000508;  wr_data_rom[ 1121]='h00000000;
    rd_cycle[ 1122] = 1'b1;  wr_cycle[ 1122] = 1'b0;  addr_rom[ 1122]='h000001e8;  wr_data_rom[ 1122]='h00000000;
    rd_cycle[ 1123] = 1'b0;  wr_cycle[ 1123] = 1'b1;  addr_rom[ 1123]='h000007fc;  wr_data_rom[ 1123]='h0000007e;
    rd_cycle[ 1124] = 1'b0;  wr_cycle[ 1124] = 1'b1;  addr_rom[ 1124]='h000005ec;  wr_data_rom[ 1124]='h00000313;
    rd_cycle[ 1125] = 1'b0;  wr_cycle[ 1125] = 1'b1;  addr_rom[ 1125]='h00000784;  wr_data_rom[ 1125]='h000001c8;
    rd_cycle[ 1126] = 1'b1;  wr_cycle[ 1126] = 1'b0;  addr_rom[ 1126]='h00000700;  wr_data_rom[ 1126]='h00000000;
    rd_cycle[ 1127] = 1'b0;  wr_cycle[ 1127] = 1'b1;  addr_rom[ 1127]='h00000004;  wr_data_rom[ 1127]='h00000236;
    rd_cycle[ 1128] = 1'b1;  wr_cycle[ 1128] = 1'b0;  addr_rom[ 1128]='h00000224;  wr_data_rom[ 1128]='h00000000;
    rd_cycle[ 1129] = 1'b1;  wr_cycle[ 1129] = 1'b0;  addr_rom[ 1129]='h000006a4;  wr_data_rom[ 1129]='h00000000;
    rd_cycle[ 1130] = 1'b1;  wr_cycle[ 1130] = 1'b0;  addr_rom[ 1130]='h00000244;  wr_data_rom[ 1130]='h00000000;
    rd_cycle[ 1131] = 1'b0;  wr_cycle[ 1131] = 1'b1;  addr_rom[ 1131]='h00000098;  wr_data_rom[ 1131]='h000002af;
    rd_cycle[ 1132] = 1'b1;  wr_cycle[ 1132] = 1'b0;  addr_rom[ 1132]='h000001b0;  wr_data_rom[ 1132]='h00000000;
    rd_cycle[ 1133] = 1'b0;  wr_cycle[ 1133] = 1'b1;  addr_rom[ 1133]='h0000033c;  wr_data_rom[ 1133]='h00000150;
    rd_cycle[ 1134] = 1'b1;  wr_cycle[ 1134] = 1'b0;  addr_rom[ 1134]='h0000030c;  wr_data_rom[ 1134]='h00000000;
    rd_cycle[ 1135] = 1'b0;  wr_cycle[ 1135] = 1'b1;  addr_rom[ 1135]='h00000650;  wr_data_rom[ 1135]='h00000618;
    rd_cycle[ 1136] = 1'b0;  wr_cycle[ 1136] = 1'b1;  addr_rom[ 1136]='h00000268;  wr_data_rom[ 1136]='h00000290;
    rd_cycle[ 1137] = 1'b1;  wr_cycle[ 1137] = 1'b0;  addr_rom[ 1137]='h00000658;  wr_data_rom[ 1137]='h00000000;
    rd_cycle[ 1138] = 1'b0;  wr_cycle[ 1138] = 1'b1;  addr_rom[ 1138]='h00000610;  wr_data_rom[ 1138]='h00000755;
    rd_cycle[ 1139] = 1'b1;  wr_cycle[ 1139] = 1'b0;  addr_rom[ 1139]='h000005b4;  wr_data_rom[ 1139]='h00000000;
    rd_cycle[ 1140] = 1'b1;  wr_cycle[ 1140] = 1'b0;  addr_rom[ 1140]='h00000428;  wr_data_rom[ 1140]='h00000000;
    rd_cycle[ 1141] = 1'b0;  wr_cycle[ 1141] = 1'b1;  addr_rom[ 1141]='h000007f4;  wr_data_rom[ 1141]='h0000002a;
    rd_cycle[ 1142] = 1'b0;  wr_cycle[ 1142] = 1'b1;  addr_rom[ 1142]='h00000688;  wr_data_rom[ 1142]='h00000225;
    rd_cycle[ 1143] = 1'b0;  wr_cycle[ 1143] = 1'b1;  addr_rom[ 1143]='h00000584;  wr_data_rom[ 1143]='h00000301;
    rd_cycle[ 1144] = 1'b1;  wr_cycle[ 1144] = 1'b0;  addr_rom[ 1144]='h000004c8;  wr_data_rom[ 1144]='h00000000;
    rd_cycle[ 1145] = 1'b1;  wr_cycle[ 1145] = 1'b0;  addr_rom[ 1145]='h00000738;  wr_data_rom[ 1145]='h00000000;
    rd_cycle[ 1146] = 1'b1;  wr_cycle[ 1146] = 1'b0;  addr_rom[ 1146]='h0000061c;  wr_data_rom[ 1146]='h00000000;
    rd_cycle[ 1147] = 1'b1;  wr_cycle[ 1147] = 1'b0;  addr_rom[ 1147]='h00000128;  wr_data_rom[ 1147]='h00000000;
    rd_cycle[ 1148] = 1'b1;  wr_cycle[ 1148] = 1'b0;  addr_rom[ 1148]='h00000310;  wr_data_rom[ 1148]='h00000000;
    rd_cycle[ 1149] = 1'b0;  wr_cycle[ 1149] = 1'b1;  addr_rom[ 1149]='h00000548;  wr_data_rom[ 1149]='h0000003f;
    rd_cycle[ 1150] = 1'b0;  wr_cycle[ 1150] = 1'b1;  addr_rom[ 1150]='h000002e0;  wr_data_rom[ 1150]='h000000ba;
    rd_cycle[ 1151] = 1'b1;  wr_cycle[ 1151] = 1'b0;  addr_rom[ 1151]='h0000010c;  wr_data_rom[ 1151]='h00000000;
    rd_cycle[ 1152] = 1'b1;  wr_cycle[ 1152] = 1'b0;  addr_rom[ 1152]='h000004f4;  wr_data_rom[ 1152]='h00000000;
    rd_cycle[ 1153] = 1'b0;  wr_cycle[ 1153] = 1'b1;  addr_rom[ 1153]='h00000774;  wr_data_rom[ 1153]='h000005fd;
    rd_cycle[ 1154] = 1'b0;  wr_cycle[ 1154] = 1'b1;  addr_rom[ 1154]='h000003e8;  wr_data_rom[ 1154]='h00000741;
    rd_cycle[ 1155] = 1'b1;  wr_cycle[ 1155] = 1'b0;  addr_rom[ 1155]='h00000688;  wr_data_rom[ 1155]='h00000000;
    rd_cycle[ 1156] = 1'b0;  wr_cycle[ 1156] = 1'b1;  addr_rom[ 1156]='h00000164;  wr_data_rom[ 1156]='h0000044e;
    rd_cycle[ 1157] = 1'b0;  wr_cycle[ 1157] = 1'b1;  addr_rom[ 1157]='h000001d0;  wr_data_rom[ 1157]='h00000200;
    rd_cycle[ 1158] = 1'b1;  wr_cycle[ 1158] = 1'b0;  addr_rom[ 1158]='h000003f0;  wr_data_rom[ 1158]='h00000000;
    rd_cycle[ 1159] = 1'b1;  wr_cycle[ 1159] = 1'b0;  addr_rom[ 1159]='h00000274;  wr_data_rom[ 1159]='h00000000;
    rd_cycle[ 1160] = 1'b1;  wr_cycle[ 1160] = 1'b0;  addr_rom[ 1160]='h00000308;  wr_data_rom[ 1160]='h00000000;
    rd_cycle[ 1161] = 1'b1;  wr_cycle[ 1161] = 1'b0;  addr_rom[ 1161]='h000003ec;  wr_data_rom[ 1161]='h00000000;
    rd_cycle[ 1162] = 1'b0;  wr_cycle[ 1162] = 1'b1;  addr_rom[ 1162]='h00000154;  wr_data_rom[ 1162]='h00000084;
    rd_cycle[ 1163] = 1'b0;  wr_cycle[ 1163] = 1'b1;  addr_rom[ 1163]='h00000470;  wr_data_rom[ 1163]='h000006d9;
    rd_cycle[ 1164] = 1'b0;  wr_cycle[ 1164] = 1'b1;  addr_rom[ 1164]='h00000120;  wr_data_rom[ 1164]='h000002e1;
    rd_cycle[ 1165] = 1'b0;  wr_cycle[ 1165] = 1'b1;  addr_rom[ 1165]='h000000fc;  wr_data_rom[ 1165]='h00000741;
    rd_cycle[ 1166] = 1'b1;  wr_cycle[ 1166] = 1'b0;  addr_rom[ 1166]='h000003c8;  wr_data_rom[ 1166]='h00000000;
    rd_cycle[ 1167] = 1'b0;  wr_cycle[ 1167] = 1'b1;  addr_rom[ 1167]='h0000014c;  wr_data_rom[ 1167]='h0000060d;
    rd_cycle[ 1168] = 1'b1;  wr_cycle[ 1168] = 1'b0;  addr_rom[ 1168]='h000000c0;  wr_data_rom[ 1168]='h00000000;
    rd_cycle[ 1169] = 1'b0;  wr_cycle[ 1169] = 1'b1;  addr_rom[ 1169]='h00000218;  wr_data_rom[ 1169]='h0000022c;
    rd_cycle[ 1170] = 1'b0;  wr_cycle[ 1170] = 1'b1;  addr_rom[ 1170]='h000007e0;  wr_data_rom[ 1170]='h000002d6;
    rd_cycle[ 1171] = 1'b1;  wr_cycle[ 1171] = 1'b0;  addr_rom[ 1171]='h000005ec;  wr_data_rom[ 1171]='h00000000;
    rd_cycle[ 1172] = 1'b1;  wr_cycle[ 1172] = 1'b0;  addr_rom[ 1172]='h000001d0;  wr_data_rom[ 1172]='h00000000;
    rd_cycle[ 1173] = 1'b0;  wr_cycle[ 1173] = 1'b1;  addr_rom[ 1173]='h0000008c;  wr_data_rom[ 1173]='h000005d0;
    rd_cycle[ 1174] = 1'b0;  wr_cycle[ 1174] = 1'b1;  addr_rom[ 1174]='h000002ec;  wr_data_rom[ 1174]='h00000483;
    rd_cycle[ 1175] = 1'b0;  wr_cycle[ 1175] = 1'b1;  addr_rom[ 1175]='h00000560;  wr_data_rom[ 1175]='h0000019e;
    rd_cycle[ 1176] = 1'b1;  wr_cycle[ 1176] = 1'b0;  addr_rom[ 1176]='h000003f8;  wr_data_rom[ 1176]='h00000000;
    rd_cycle[ 1177] = 1'b0;  wr_cycle[ 1177] = 1'b1;  addr_rom[ 1177]='h00000534;  wr_data_rom[ 1177]='h00000166;
    rd_cycle[ 1178] = 1'b0;  wr_cycle[ 1178] = 1'b1;  addr_rom[ 1178]='h0000003c;  wr_data_rom[ 1178]='h0000022f;
    rd_cycle[ 1179] = 1'b1;  wr_cycle[ 1179] = 1'b0;  addr_rom[ 1179]='h000006c4;  wr_data_rom[ 1179]='h00000000;
    rd_cycle[ 1180] = 1'b1;  wr_cycle[ 1180] = 1'b0;  addr_rom[ 1180]='h000005fc;  wr_data_rom[ 1180]='h00000000;
    rd_cycle[ 1181] = 1'b1;  wr_cycle[ 1181] = 1'b0;  addr_rom[ 1181]='h000005a4;  wr_data_rom[ 1181]='h00000000;
    rd_cycle[ 1182] = 1'b0;  wr_cycle[ 1182] = 1'b1;  addr_rom[ 1182]='h000006a0;  wr_data_rom[ 1182]='h000002d3;
    rd_cycle[ 1183] = 1'b1;  wr_cycle[ 1183] = 1'b0;  addr_rom[ 1183]='h00000488;  wr_data_rom[ 1183]='h00000000;
    rd_cycle[ 1184] = 1'b0;  wr_cycle[ 1184] = 1'b1;  addr_rom[ 1184]='h00000068;  wr_data_rom[ 1184]='h00000701;
    rd_cycle[ 1185] = 1'b0;  wr_cycle[ 1185] = 1'b1;  addr_rom[ 1185]='h000000b4;  wr_data_rom[ 1185]='h0000011a;
    rd_cycle[ 1186] = 1'b0;  wr_cycle[ 1186] = 1'b1;  addr_rom[ 1186]='h00000638;  wr_data_rom[ 1186]='h000002cc;
    rd_cycle[ 1187] = 1'b0;  wr_cycle[ 1187] = 1'b1;  addr_rom[ 1187]='h000003dc;  wr_data_rom[ 1187]='h0000007b;
    rd_cycle[ 1188] = 1'b0;  wr_cycle[ 1188] = 1'b1;  addr_rom[ 1188]='h00000548;  wr_data_rom[ 1188]='h000006c6;
    rd_cycle[ 1189] = 1'b1;  wr_cycle[ 1189] = 1'b0;  addr_rom[ 1189]='h0000013c;  wr_data_rom[ 1189]='h00000000;
    rd_cycle[ 1190] = 1'b0;  wr_cycle[ 1190] = 1'b1;  addr_rom[ 1190]='h000002e4;  wr_data_rom[ 1190]='h000005cf;
    rd_cycle[ 1191] = 1'b1;  wr_cycle[ 1191] = 1'b0;  addr_rom[ 1191]='h00000124;  wr_data_rom[ 1191]='h00000000;
    rd_cycle[ 1192] = 1'b0;  wr_cycle[ 1192] = 1'b1;  addr_rom[ 1192]='h0000036c;  wr_data_rom[ 1192]='h00000644;
    rd_cycle[ 1193] = 1'b1;  wr_cycle[ 1193] = 1'b0;  addr_rom[ 1193]='h000000a0;  wr_data_rom[ 1193]='h00000000;
    rd_cycle[ 1194] = 1'b1;  wr_cycle[ 1194] = 1'b0;  addr_rom[ 1194]='h00000230;  wr_data_rom[ 1194]='h00000000;
    rd_cycle[ 1195] = 1'b1;  wr_cycle[ 1195] = 1'b0;  addr_rom[ 1195]='h00000594;  wr_data_rom[ 1195]='h00000000;
    rd_cycle[ 1196] = 1'b1;  wr_cycle[ 1196] = 1'b0;  addr_rom[ 1196]='h00000324;  wr_data_rom[ 1196]='h00000000;
    rd_cycle[ 1197] = 1'b1;  wr_cycle[ 1197] = 1'b0;  addr_rom[ 1197]='h000005a4;  wr_data_rom[ 1197]='h00000000;
    rd_cycle[ 1198] = 1'b0;  wr_cycle[ 1198] = 1'b1;  addr_rom[ 1198]='h00000014;  wr_data_rom[ 1198]='h000006d7;
    rd_cycle[ 1199] = 1'b1;  wr_cycle[ 1199] = 1'b0;  addr_rom[ 1199]='h000002f0;  wr_data_rom[ 1199]='h00000000;
    rd_cycle[ 1200] = 1'b0;  wr_cycle[ 1200] = 1'b1;  addr_rom[ 1200]='h0000031c;  wr_data_rom[ 1200]='h00000237;
    rd_cycle[ 1201] = 1'b1;  wr_cycle[ 1201] = 1'b0;  addr_rom[ 1201]='h00000378;  wr_data_rom[ 1201]='h00000000;
    rd_cycle[ 1202] = 1'b0;  wr_cycle[ 1202] = 1'b1;  addr_rom[ 1202]='h000002e0;  wr_data_rom[ 1202]='h000001a6;
    rd_cycle[ 1203] = 1'b1;  wr_cycle[ 1203] = 1'b0;  addr_rom[ 1203]='h00000110;  wr_data_rom[ 1203]='h00000000;
    rd_cycle[ 1204] = 1'b1;  wr_cycle[ 1204] = 1'b0;  addr_rom[ 1204]='h000005fc;  wr_data_rom[ 1204]='h00000000;
    rd_cycle[ 1205] = 1'b0;  wr_cycle[ 1205] = 1'b1;  addr_rom[ 1205]='h0000075c;  wr_data_rom[ 1205]='h00000556;
    rd_cycle[ 1206] = 1'b0;  wr_cycle[ 1206] = 1'b1;  addr_rom[ 1206]='h000004a0;  wr_data_rom[ 1206]='h000006ec;
    rd_cycle[ 1207] = 1'b0;  wr_cycle[ 1207] = 1'b1;  addr_rom[ 1207]='h00000034;  wr_data_rom[ 1207]='h000007f1;
    rd_cycle[ 1208] = 1'b1;  wr_cycle[ 1208] = 1'b0;  addr_rom[ 1208]='h000000b4;  wr_data_rom[ 1208]='h00000000;
    rd_cycle[ 1209] = 1'b0;  wr_cycle[ 1209] = 1'b1;  addr_rom[ 1209]='h00000734;  wr_data_rom[ 1209]='h00000669;
    rd_cycle[ 1210] = 1'b1;  wr_cycle[ 1210] = 1'b0;  addr_rom[ 1210]='h00000204;  wr_data_rom[ 1210]='h00000000;
    rd_cycle[ 1211] = 1'b0;  wr_cycle[ 1211] = 1'b1;  addr_rom[ 1211]='h00000358;  wr_data_rom[ 1211]='h0000031d;
    rd_cycle[ 1212] = 1'b1;  wr_cycle[ 1212] = 1'b0;  addr_rom[ 1212]='h000003a0;  wr_data_rom[ 1212]='h00000000;
    rd_cycle[ 1213] = 1'b0;  wr_cycle[ 1213] = 1'b1;  addr_rom[ 1213]='h0000034c;  wr_data_rom[ 1213]='h00000143;
    rd_cycle[ 1214] = 1'b1;  wr_cycle[ 1214] = 1'b0;  addr_rom[ 1214]='h0000070c;  wr_data_rom[ 1214]='h00000000;
    rd_cycle[ 1215] = 1'b1;  wr_cycle[ 1215] = 1'b0;  addr_rom[ 1215]='h00000660;  wr_data_rom[ 1215]='h00000000;
    rd_cycle[ 1216] = 1'b0;  wr_cycle[ 1216] = 1'b1;  addr_rom[ 1216]='h0000008c;  wr_data_rom[ 1216]='h000003bb;
    rd_cycle[ 1217] = 1'b0;  wr_cycle[ 1217] = 1'b1;  addr_rom[ 1217]='h000000b8;  wr_data_rom[ 1217]='h00000012;
    rd_cycle[ 1218] = 1'b0;  wr_cycle[ 1218] = 1'b1;  addr_rom[ 1218]='h00000044;  wr_data_rom[ 1218]='h00000772;
    rd_cycle[ 1219] = 1'b0;  wr_cycle[ 1219] = 1'b1;  addr_rom[ 1219]='h000002a8;  wr_data_rom[ 1219]='h0000005d;
    rd_cycle[ 1220] = 1'b1;  wr_cycle[ 1220] = 1'b0;  addr_rom[ 1220]='h00000180;  wr_data_rom[ 1220]='h00000000;
    rd_cycle[ 1221] = 1'b0;  wr_cycle[ 1221] = 1'b1;  addr_rom[ 1221]='h0000024c;  wr_data_rom[ 1221]='h000000e2;
    rd_cycle[ 1222] = 1'b1;  wr_cycle[ 1222] = 1'b0;  addr_rom[ 1222]='h00000564;  wr_data_rom[ 1222]='h00000000;
    rd_cycle[ 1223] = 1'b1;  wr_cycle[ 1223] = 1'b0;  addr_rom[ 1223]='h00000684;  wr_data_rom[ 1223]='h00000000;
    rd_cycle[ 1224] = 1'b0;  wr_cycle[ 1224] = 1'b1;  addr_rom[ 1224]='h00000068;  wr_data_rom[ 1224]='h00000005;
    rd_cycle[ 1225] = 1'b1;  wr_cycle[ 1225] = 1'b0;  addr_rom[ 1225]='h0000002c;  wr_data_rom[ 1225]='h00000000;
    rd_cycle[ 1226] = 1'b0;  wr_cycle[ 1226] = 1'b1;  addr_rom[ 1226]='h00000244;  wr_data_rom[ 1226]='h0000023a;
    rd_cycle[ 1227] = 1'b1;  wr_cycle[ 1227] = 1'b0;  addr_rom[ 1227]='h0000074c;  wr_data_rom[ 1227]='h00000000;
    rd_cycle[ 1228] = 1'b0;  wr_cycle[ 1228] = 1'b1;  addr_rom[ 1228]='h000000e0;  wr_data_rom[ 1228]='h0000055f;
    rd_cycle[ 1229] = 1'b0;  wr_cycle[ 1229] = 1'b1;  addr_rom[ 1229]='h00000508;  wr_data_rom[ 1229]='h000006a6;
    rd_cycle[ 1230] = 1'b0;  wr_cycle[ 1230] = 1'b1;  addr_rom[ 1230]='h000001fc;  wr_data_rom[ 1230]='h00000062;
    rd_cycle[ 1231] = 1'b1;  wr_cycle[ 1231] = 1'b0;  addr_rom[ 1231]='h00000200;  wr_data_rom[ 1231]='h00000000;
    rd_cycle[ 1232] = 1'b1;  wr_cycle[ 1232] = 1'b0;  addr_rom[ 1232]='h0000031c;  wr_data_rom[ 1232]='h00000000;
    rd_cycle[ 1233] = 1'b0;  wr_cycle[ 1233] = 1'b1;  addr_rom[ 1233]='h00000328;  wr_data_rom[ 1233]='h000000c8;
    rd_cycle[ 1234] = 1'b1;  wr_cycle[ 1234] = 1'b0;  addr_rom[ 1234]='h00000218;  wr_data_rom[ 1234]='h00000000;
    rd_cycle[ 1235] = 1'b0;  wr_cycle[ 1235] = 1'b1;  addr_rom[ 1235]='h0000043c;  wr_data_rom[ 1235]='h00000029;
    rd_cycle[ 1236] = 1'b0;  wr_cycle[ 1236] = 1'b1;  addr_rom[ 1236]='h00000780;  wr_data_rom[ 1236]='h000007ae;
    rd_cycle[ 1237] = 1'b0;  wr_cycle[ 1237] = 1'b1;  addr_rom[ 1237]='h000005c0;  wr_data_rom[ 1237]='h00000163;
    rd_cycle[ 1238] = 1'b0;  wr_cycle[ 1238] = 1'b1;  addr_rom[ 1238]='h00000250;  wr_data_rom[ 1238]='h000000ec;
    rd_cycle[ 1239] = 1'b1;  wr_cycle[ 1239] = 1'b0;  addr_rom[ 1239]='h00000640;  wr_data_rom[ 1239]='h00000000;
    rd_cycle[ 1240] = 1'b0;  wr_cycle[ 1240] = 1'b1;  addr_rom[ 1240]='h00000120;  wr_data_rom[ 1240]='h000002bb;
    rd_cycle[ 1241] = 1'b0;  wr_cycle[ 1241] = 1'b1;  addr_rom[ 1241]='h000004c8;  wr_data_rom[ 1241]='h0000020c;
    rd_cycle[ 1242] = 1'b0;  wr_cycle[ 1242] = 1'b1;  addr_rom[ 1242]='h00000798;  wr_data_rom[ 1242]='h000003a3;
    rd_cycle[ 1243] = 1'b0;  wr_cycle[ 1243] = 1'b1;  addr_rom[ 1243]='h000004d4;  wr_data_rom[ 1243]='h0000079f;
    rd_cycle[ 1244] = 1'b0;  wr_cycle[ 1244] = 1'b1;  addr_rom[ 1244]='h000005fc;  wr_data_rom[ 1244]='h000000b9;
    rd_cycle[ 1245] = 1'b0;  wr_cycle[ 1245] = 1'b1;  addr_rom[ 1245]='h00000130;  wr_data_rom[ 1245]='h00000486;
    rd_cycle[ 1246] = 1'b1;  wr_cycle[ 1246] = 1'b0;  addr_rom[ 1246]='h00000654;  wr_data_rom[ 1246]='h00000000;
    rd_cycle[ 1247] = 1'b1;  wr_cycle[ 1247] = 1'b0;  addr_rom[ 1247]='h00000460;  wr_data_rom[ 1247]='h00000000;
    rd_cycle[ 1248] = 1'b0;  wr_cycle[ 1248] = 1'b1;  addr_rom[ 1248]='h00000440;  wr_data_rom[ 1248]='h00000028;
    rd_cycle[ 1249] = 1'b0;  wr_cycle[ 1249] = 1'b1;  addr_rom[ 1249]='h0000062c;  wr_data_rom[ 1249]='h000002c9;
    rd_cycle[ 1250] = 1'b0;  wr_cycle[ 1250] = 1'b1;  addr_rom[ 1250]='h000004e8;  wr_data_rom[ 1250]='h00000447;
    rd_cycle[ 1251] = 1'b1;  wr_cycle[ 1251] = 1'b0;  addr_rom[ 1251]='h0000013c;  wr_data_rom[ 1251]='h00000000;
    rd_cycle[ 1252] = 1'b1;  wr_cycle[ 1252] = 1'b0;  addr_rom[ 1252]='h000005ac;  wr_data_rom[ 1252]='h00000000;
    rd_cycle[ 1253] = 1'b1;  wr_cycle[ 1253] = 1'b0;  addr_rom[ 1253]='h00000454;  wr_data_rom[ 1253]='h00000000;
    rd_cycle[ 1254] = 1'b1;  wr_cycle[ 1254] = 1'b0;  addr_rom[ 1254]='h00000148;  wr_data_rom[ 1254]='h00000000;
    rd_cycle[ 1255] = 1'b0;  wr_cycle[ 1255] = 1'b1;  addr_rom[ 1255]='h00000004;  wr_data_rom[ 1255]='h000001b9;
    rd_cycle[ 1256] = 1'b0;  wr_cycle[ 1256] = 1'b1;  addr_rom[ 1256]='h0000046c;  wr_data_rom[ 1256]='h0000008f;
    rd_cycle[ 1257] = 1'b0;  wr_cycle[ 1257] = 1'b1;  addr_rom[ 1257]='h000007e0;  wr_data_rom[ 1257]='h0000073a;
    rd_cycle[ 1258] = 1'b1;  wr_cycle[ 1258] = 1'b0;  addr_rom[ 1258]='h000004b8;  wr_data_rom[ 1258]='h00000000;
    rd_cycle[ 1259] = 1'b1;  wr_cycle[ 1259] = 1'b0;  addr_rom[ 1259]='h000006f0;  wr_data_rom[ 1259]='h00000000;
    rd_cycle[ 1260] = 1'b1;  wr_cycle[ 1260] = 1'b0;  addr_rom[ 1260]='h00000140;  wr_data_rom[ 1260]='h00000000;
    rd_cycle[ 1261] = 1'b0;  wr_cycle[ 1261] = 1'b1;  addr_rom[ 1261]='h000003c8;  wr_data_rom[ 1261]='h00000735;
    rd_cycle[ 1262] = 1'b1;  wr_cycle[ 1262] = 1'b0;  addr_rom[ 1262]='h000004e0;  wr_data_rom[ 1262]='h00000000;
    rd_cycle[ 1263] = 1'b0;  wr_cycle[ 1263] = 1'b1;  addr_rom[ 1263]='h000005f0;  wr_data_rom[ 1263]='h000004f5;
    rd_cycle[ 1264] = 1'b1;  wr_cycle[ 1264] = 1'b0;  addr_rom[ 1264]='h0000064c;  wr_data_rom[ 1264]='h00000000;
    rd_cycle[ 1265] = 1'b1;  wr_cycle[ 1265] = 1'b0;  addr_rom[ 1265]='h0000070c;  wr_data_rom[ 1265]='h00000000;
    rd_cycle[ 1266] = 1'b1;  wr_cycle[ 1266] = 1'b0;  addr_rom[ 1266]='h0000004c;  wr_data_rom[ 1266]='h00000000;
    rd_cycle[ 1267] = 1'b1;  wr_cycle[ 1267] = 1'b0;  addr_rom[ 1267]='h000002a0;  wr_data_rom[ 1267]='h00000000;
    rd_cycle[ 1268] = 1'b0;  wr_cycle[ 1268] = 1'b1;  addr_rom[ 1268]='h000000ac;  wr_data_rom[ 1268]='h0000041a;
    rd_cycle[ 1269] = 1'b1;  wr_cycle[ 1269] = 1'b0;  addr_rom[ 1269]='h00000660;  wr_data_rom[ 1269]='h00000000;
    rd_cycle[ 1270] = 1'b0;  wr_cycle[ 1270] = 1'b1;  addr_rom[ 1270]='h00000204;  wr_data_rom[ 1270]='h0000020e;
    rd_cycle[ 1271] = 1'b0;  wr_cycle[ 1271] = 1'b1;  addr_rom[ 1271]='h000002c0;  wr_data_rom[ 1271]='h00000621;
    rd_cycle[ 1272] = 1'b1;  wr_cycle[ 1272] = 1'b0;  addr_rom[ 1272]='h00000644;  wr_data_rom[ 1272]='h00000000;
    rd_cycle[ 1273] = 1'b1;  wr_cycle[ 1273] = 1'b0;  addr_rom[ 1273]='h000006ec;  wr_data_rom[ 1273]='h00000000;
    rd_cycle[ 1274] = 1'b1;  wr_cycle[ 1274] = 1'b0;  addr_rom[ 1274]='h0000059c;  wr_data_rom[ 1274]='h00000000;
    rd_cycle[ 1275] = 1'b0;  wr_cycle[ 1275] = 1'b1;  addr_rom[ 1275]='h000001f8;  wr_data_rom[ 1275]='h000004eb;
    rd_cycle[ 1276] = 1'b1;  wr_cycle[ 1276] = 1'b0;  addr_rom[ 1276]='h000006f8;  wr_data_rom[ 1276]='h00000000;
    rd_cycle[ 1277] = 1'b0;  wr_cycle[ 1277] = 1'b1;  addr_rom[ 1277]='h00000004;  wr_data_rom[ 1277]='h00000450;
    rd_cycle[ 1278] = 1'b1;  wr_cycle[ 1278] = 1'b0;  addr_rom[ 1278]='h00000784;  wr_data_rom[ 1278]='h00000000;
    rd_cycle[ 1279] = 1'b0;  wr_cycle[ 1279] = 1'b1;  addr_rom[ 1279]='h0000010c;  wr_data_rom[ 1279]='h00000083;
    rd_cycle[ 1280] = 1'b1;  wr_cycle[ 1280] = 1'b0;  addr_rom[ 1280]='h000006d0;  wr_data_rom[ 1280]='h00000000;
    rd_cycle[ 1281] = 1'b1;  wr_cycle[ 1281] = 1'b0;  addr_rom[ 1281]='h000006ec;  wr_data_rom[ 1281]='h00000000;
    rd_cycle[ 1282] = 1'b1;  wr_cycle[ 1282] = 1'b0;  addr_rom[ 1282]='h0000002c;  wr_data_rom[ 1282]='h00000000;
    rd_cycle[ 1283] = 1'b1;  wr_cycle[ 1283] = 1'b0;  addr_rom[ 1283]='h0000072c;  wr_data_rom[ 1283]='h00000000;
    rd_cycle[ 1284] = 1'b1;  wr_cycle[ 1284] = 1'b0;  addr_rom[ 1284]='h0000034c;  wr_data_rom[ 1284]='h00000000;
    rd_cycle[ 1285] = 1'b0;  wr_cycle[ 1285] = 1'b1;  addr_rom[ 1285]='h00000090;  wr_data_rom[ 1285]='h000006b2;
    rd_cycle[ 1286] = 1'b1;  wr_cycle[ 1286] = 1'b0;  addr_rom[ 1286]='h000004a4;  wr_data_rom[ 1286]='h00000000;
    rd_cycle[ 1287] = 1'b1;  wr_cycle[ 1287] = 1'b0;  addr_rom[ 1287]='h00000594;  wr_data_rom[ 1287]='h00000000;
    rd_cycle[ 1288] = 1'b1;  wr_cycle[ 1288] = 1'b0;  addr_rom[ 1288]='h000003c0;  wr_data_rom[ 1288]='h00000000;
    rd_cycle[ 1289] = 1'b0;  wr_cycle[ 1289] = 1'b1;  addr_rom[ 1289]='h000000e8;  wr_data_rom[ 1289]='h000001aa;
    rd_cycle[ 1290] = 1'b1;  wr_cycle[ 1290] = 1'b0;  addr_rom[ 1290]='h000002a0;  wr_data_rom[ 1290]='h00000000;
    rd_cycle[ 1291] = 1'b1;  wr_cycle[ 1291] = 1'b0;  addr_rom[ 1291]='h000007c8;  wr_data_rom[ 1291]='h00000000;
    rd_cycle[ 1292] = 1'b0;  wr_cycle[ 1292] = 1'b1;  addr_rom[ 1292]='h000001a8;  wr_data_rom[ 1292]='h000004eb;
    rd_cycle[ 1293] = 1'b1;  wr_cycle[ 1293] = 1'b0;  addr_rom[ 1293]='h00000238;  wr_data_rom[ 1293]='h00000000;
    rd_cycle[ 1294] = 1'b0;  wr_cycle[ 1294] = 1'b1;  addr_rom[ 1294]='h00000440;  wr_data_rom[ 1294]='h000004c3;
    rd_cycle[ 1295] = 1'b0;  wr_cycle[ 1295] = 1'b1;  addr_rom[ 1295]='h000002c4;  wr_data_rom[ 1295]='h000005d4;
    rd_cycle[ 1296] = 1'b0;  wr_cycle[ 1296] = 1'b1;  addr_rom[ 1296]='h000001c4;  wr_data_rom[ 1296]='h0000064d;
    rd_cycle[ 1297] = 1'b0;  wr_cycle[ 1297] = 1'b1;  addr_rom[ 1297]='h0000002c;  wr_data_rom[ 1297]='h0000039d;
    rd_cycle[ 1298] = 1'b0;  wr_cycle[ 1298] = 1'b1;  addr_rom[ 1298]='h00000414;  wr_data_rom[ 1298]='h000004d5;
    rd_cycle[ 1299] = 1'b1;  wr_cycle[ 1299] = 1'b0;  addr_rom[ 1299]='h00000670;  wr_data_rom[ 1299]='h00000000;
    rd_cycle[ 1300] = 1'b1;  wr_cycle[ 1300] = 1'b0;  addr_rom[ 1300]='h0000024c;  wr_data_rom[ 1300]='h00000000;
    rd_cycle[ 1301] = 1'b0;  wr_cycle[ 1301] = 1'b1;  addr_rom[ 1301]='h000007b8;  wr_data_rom[ 1301]='h00000255;
    rd_cycle[ 1302] = 1'b0;  wr_cycle[ 1302] = 1'b1;  addr_rom[ 1302]='h00000080;  wr_data_rom[ 1302]='h000004be;
    rd_cycle[ 1303] = 1'b0;  wr_cycle[ 1303] = 1'b1;  addr_rom[ 1303]='h00000280;  wr_data_rom[ 1303]='h000002a6;
    rd_cycle[ 1304] = 1'b1;  wr_cycle[ 1304] = 1'b0;  addr_rom[ 1304]='h00000728;  wr_data_rom[ 1304]='h00000000;
    rd_cycle[ 1305] = 1'b1;  wr_cycle[ 1305] = 1'b0;  addr_rom[ 1305]='h00000434;  wr_data_rom[ 1305]='h00000000;
    rd_cycle[ 1306] = 1'b0;  wr_cycle[ 1306] = 1'b1;  addr_rom[ 1306]='h000006c0;  wr_data_rom[ 1306]='h000007b0;
    rd_cycle[ 1307] = 1'b0;  wr_cycle[ 1307] = 1'b1;  addr_rom[ 1307]='h00000484;  wr_data_rom[ 1307]='h0000065d;
    rd_cycle[ 1308] = 1'b1;  wr_cycle[ 1308] = 1'b0;  addr_rom[ 1308]='h0000036c;  wr_data_rom[ 1308]='h00000000;
    rd_cycle[ 1309] = 1'b0;  wr_cycle[ 1309] = 1'b1;  addr_rom[ 1309]='h0000028c;  wr_data_rom[ 1309]='h0000022e;
    rd_cycle[ 1310] = 1'b1;  wr_cycle[ 1310] = 1'b0;  addr_rom[ 1310]='h0000032c;  wr_data_rom[ 1310]='h00000000;
    rd_cycle[ 1311] = 1'b1;  wr_cycle[ 1311] = 1'b0;  addr_rom[ 1311]='h00000630;  wr_data_rom[ 1311]='h00000000;
    rd_cycle[ 1312] = 1'b1;  wr_cycle[ 1312] = 1'b0;  addr_rom[ 1312]='h000006f0;  wr_data_rom[ 1312]='h00000000;
    rd_cycle[ 1313] = 1'b0;  wr_cycle[ 1313] = 1'b1;  addr_rom[ 1313]='h0000064c;  wr_data_rom[ 1313]='h0000026f;
    rd_cycle[ 1314] = 1'b0;  wr_cycle[ 1314] = 1'b1;  addr_rom[ 1314]='h000004fc;  wr_data_rom[ 1314]='h00000342;
    rd_cycle[ 1315] = 1'b1;  wr_cycle[ 1315] = 1'b0;  addr_rom[ 1315]='h000005a8;  wr_data_rom[ 1315]='h00000000;
    rd_cycle[ 1316] = 1'b0;  wr_cycle[ 1316] = 1'b1;  addr_rom[ 1316]='h000003b4;  wr_data_rom[ 1316]='h0000001d;
    rd_cycle[ 1317] = 1'b0;  wr_cycle[ 1317] = 1'b1;  addr_rom[ 1317]='h0000053c;  wr_data_rom[ 1317]='h000003dd;
    rd_cycle[ 1318] = 1'b0;  wr_cycle[ 1318] = 1'b1;  addr_rom[ 1318]='h00000350;  wr_data_rom[ 1318]='h000006e7;
    rd_cycle[ 1319] = 1'b1;  wr_cycle[ 1319] = 1'b0;  addr_rom[ 1319]='h00000784;  wr_data_rom[ 1319]='h00000000;
    rd_cycle[ 1320] = 1'b0;  wr_cycle[ 1320] = 1'b1;  addr_rom[ 1320]='h000007b4;  wr_data_rom[ 1320]='h000005ad;
    rd_cycle[ 1321] = 1'b1;  wr_cycle[ 1321] = 1'b0;  addr_rom[ 1321]='h00000688;  wr_data_rom[ 1321]='h00000000;
    rd_cycle[ 1322] = 1'b0;  wr_cycle[ 1322] = 1'b1;  addr_rom[ 1322]='h00000270;  wr_data_rom[ 1322]='h000001f7;
    rd_cycle[ 1323] = 1'b1;  wr_cycle[ 1323] = 1'b0;  addr_rom[ 1323]='h00000068;  wr_data_rom[ 1323]='h00000000;
    rd_cycle[ 1324] = 1'b1;  wr_cycle[ 1324] = 1'b0;  addr_rom[ 1324]='h000006bc;  wr_data_rom[ 1324]='h00000000;
    rd_cycle[ 1325] = 1'b1;  wr_cycle[ 1325] = 1'b0;  addr_rom[ 1325]='h000007f4;  wr_data_rom[ 1325]='h00000000;
    rd_cycle[ 1326] = 1'b0;  wr_cycle[ 1326] = 1'b1;  addr_rom[ 1326]='h00000348;  wr_data_rom[ 1326]='h0000070a;
    rd_cycle[ 1327] = 1'b1;  wr_cycle[ 1327] = 1'b0;  addr_rom[ 1327]='h000004b0;  wr_data_rom[ 1327]='h00000000;
    rd_cycle[ 1328] = 1'b0;  wr_cycle[ 1328] = 1'b1;  addr_rom[ 1328]='h00000124;  wr_data_rom[ 1328]='h000001fb;
    rd_cycle[ 1329] = 1'b0;  wr_cycle[ 1329] = 1'b1;  addr_rom[ 1329]='h000007fc;  wr_data_rom[ 1329]='h00000694;
    rd_cycle[ 1330] = 1'b1;  wr_cycle[ 1330] = 1'b0;  addr_rom[ 1330]='h0000031c;  wr_data_rom[ 1330]='h00000000;
    rd_cycle[ 1331] = 1'b0;  wr_cycle[ 1331] = 1'b1;  addr_rom[ 1331]='h00000108;  wr_data_rom[ 1331]='h00000761;
    rd_cycle[ 1332] = 1'b0;  wr_cycle[ 1332] = 1'b1;  addr_rom[ 1332]='h0000074c;  wr_data_rom[ 1332]='h000005b8;
    rd_cycle[ 1333] = 1'b1;  wr_cycle[ 1333] = 1'b0;  addr_rom[ 1333]='h00000374;  wr_data_rom[ 1333]='h00000000;
    rd_cycle[ 1334] = 1'b0;  wr_cycle[ 1334] = 1'b1;  addr_rom[ 1334]='h000007f4;  wr_data_rom[ 1334]='h000007d6;
    rd_cycle[ 1335] = 1'b1;  wr_cycle[ 1335] = 1'b0;  addr_rom[ 1335]='h000000bc;  wr_data_rom[ 1335]='h00000000;
    rd_cycle[ 1336] = 1'b1;  wr_cycle[ 1336] = 1'b0;  addr_rom[ 1336]='h0000007c;  wr_data_rom[ 1336]='h00000000;
    rd_cycle[ 1337] = 1'b1;  wr_cycle[ 1337] = 1'b0;  addr_rom[ 1337]='h0000044c;  wr_data_rom[ 1337]='h00000000;
    rd_cycle[ 1338] = 1'b1;  wr_cycle[ 1338] = 1'b0;  addr_rom[ 1338]='h00000130;  wr_data_rom[ 1338]='h00000000;
    rd_cycle[ 1339] = 1'b1;  wr_cycle[ 1339] = 1'b0;  addr_rom[ 1339]='h00000570;  wr_data_rom[ 1339]='h00000000;
    rd_cycle[ 1340] = 1'b0;  wr_cycle[ 1340] = 1'b1;  addr_rom[ 1340]='h00000490;  wr_data_rom[ 1340]='h00000170;
    rd_cycle[ 1341] = 1'b0;  wr_cycle[ 1341] = 1'b1;  addr_rom[ 1341]='h0000074c;  wr_data_rom[ 1341]='h00000106;
    rd_cycle[ 1342] = 1'b1;  wr_cycle[ 1342] = 1'b0;  addr_rom[ 1342]='h00000390;  wr_data_rom[ 1342]='h00000000;
    rd_cycle[ 1343] = 1'b0;  wr_cycle[ 1343] = 1'b1;  addr_rom[ 1343]='h000004dc;  wr_data_rom[ 1343]='h00000693;
    rd_cycle[ 1344] = 1'b1;  wr_cycle[ 1344] = 1'b0;  addr_rom[ 1344]='h000004c8;  wr_data_rom[ 1344]='h00000000;
    rd_cycle[ 1345] = 1'b1;  wr_cycle[ 1345] = 1'b0;  addr_rom[ 1345]='h0000056c;  wr_data_rom[ 1345]='h00000000;
    rd_cycle[ 1346] = 1'b0;  wr_cycle[ 1346] = 1'b1;  addr_rom[ 1346]='h0000078c;  wr_data_rom[ 1346]='h00000479;
    rd_cycle[ 1347] = 1'b1;  wr_cycle[ 1347] = 1'b0;  addr_rom[ 1347]='h00000374;  wr_data_rom[ 1347]='h00000000;
    rd_cycle[ 1348] = 1'b0;  wr_cycle[ 1348] = 1'b1;  addr_rom[ 1348]='h000007c8;  wr_data_rom[ 1348]='h0000079e;
    rd_cycle[ 1349] = 1'b1;  wr_cycle[ 1349] = 1'b0;  addr_rom[ 1349]='h00000234;  wr_data_rom[ 1349]='h00000000;
    rd_cycle[ 1350] = 1'b0;  wr_cycle[ 1350] = 1'b1;  addr_rom[ 1350]='h000004a4;  wr_data_rom[ 1350]='h00000363;
    rd_cycle[ 1351] = 1'b0;  wr_cycle[ 1351] = 1'b1;  addr_rom[ 1351]='h000000f8;  wr_data_rom[ 1351]='h000000e4;
    rd_cycle[ 1352] = 1'b1;  wr_cycle[ 1352] = 1'b0;  addr_rom[ 1352]='h00000318;  wr_data_rom[ 1352]='h00000000;
    rd_cycle[ 1353] = 1'b1;  wr_cycle[ 1353] = 1'b0;  addr_rom[ 1353]='h000002f4;  wr_data_rom[ 1353]='h00000000;
    rd_cycle[ 1354] = 1'b0;  wr_cycle[ 1354] = 1'b1;  addr_rom[ 1354]='h000006a4;  wr_data_rom[ 1354]='h000005ae;
    rd_cycle[ 1355] = 1'b1;  wr_cycle[ 1355] = 1'b0;  addr_rom[ 1355]='h000006ac;  wr_data_rom[ 1355]='h00000000;
    rd_cycle[ 1356] = 1'b1;  wr_cycle[ 1356] = 1'b0;  addr_rom[ 1356]='h0000052c;  wr_data_rom[ 1356]='h00000000;
    rd_cycle[ 1357] = 1'b0;  wr_cycle[ 1357] = 1'b1;  addr_rom[ 1357]='h000002ec;  wr_data_rom[ 1357]='h00000638;
    rd_cycle[ 1358] = 1'b1;  wr_cycle[ 1358] = 1'b0;  addr_rom[ 1358]='h000005a4;  wr_data_rom[ 1358]='h00000000;
    rd_cycle[ 1359] = 1'b0;  wr_cycle[ 1359] = 1'b1;  addr_rom[ 1359]='h00000150;  wr_data_rom[ 1359]='h000003b1;
    rd_cycle[ 1360] = 1'b1;  wr_cycle[ 1360] = 1'b0;  addr_rom[ 1360]='h00000258;  wr_data_rom[ 1360]='h00000000;
    rd_cycle[ 1361] = 1'b0;  wr_cycle[ 1361] = 1'b1;  addr_rom[ 1361]='h000007e8;  wr_data_rom[ 1361]='h00000500;
    rd_cycle[ 1362] = 1'b1;  wr_cycle[ 1362] = 1'b0;  addr_rom[ 1362]='h00000550;  wr_data_rom[ 1362]='h00000000;
    rd_cycle[ 1363] = 1'b1;  wr_cycle[ 1363] = 1'b0;  addr_rom[ 1363]='h000000c8;  wr_data_rom[ 1363]='h00000000;
    rd_cycle[ 1364] = 1'b0;  wr_cycle[ 1364] = 1'b1;  addr_rom[ 1364]='h00000034;  wr_data_rom[ 1364]='h00000386;
    rd_cycle[ 1365] = 1'b0;  wr_cycle[ 1365] = 1'b1;  addr_rom[ 1365]='h00000554;  wr_data_rom[ 1365]='h000006df;
    rd_cycle[ 1366] = 1'b0;  wr_cycle[ 1366] = 1'b1;  addr_rom[ 1366]='h000006f8;  wr_data_rom[ 1366]='h00000307;
    rd_cycle[ 1367] = 1'b1;  wr_cycle[ 1367] = 1'b0;  addr_rom[ 1367]='h00000008;  wr_data_rom[ 1367]='h00000000;
    rd_cycle[ 1368] = 1'b1;  wr_cycle[ 1368] = 1'b0;  addr_rom[ 1368]='h000000b8;  wr_data_rom[ 1368]='h00000000;
    rd_cycle[ 1369] = 1'b0;  wr_cycle[ 1369] = 1'b1;  addr_rom[ 1369]='h00000648;  wr_data_rom[ 1369]='h00000475;
    rd_cycle[ 1370] = 1'b0;  wr_cycle[ 1370] = 1'b1;  addr_rom[ 1370]='h00000544;  wr_data_rom[ 1370]='h00000542;
    rd_cycle[ 1371] = 1'b1;  wr_cycle[ 1371] = 1'b0;  addr_rom[ 1371]='h000005d8;  wr_data_rom[ 1371]='h00000000;
    rd_cycle[ 1372] = 1'b1;  wr_cycle[ 1372] = 1'b0;  addr_rom[ 1372]='h00000470;  wr_data_rom[ 1372]='h00000000;
    rd_cycle[ 1373] = 1'b1;  wr_cycle[ 1373] = 1'b0;  addr_rom[ 1373]='h000006ac;  wr_data_rom[ 1373]='h00000000;
    rd_cycle[ 1374] = 1'b1;  wr_cycle[ 1374] = 1'b0;  addr_rom[ 1374]='h00000324;  wr_data_rom[ 1374]='h00000000;
    rd_cycle[ 1375] = 1'b0;  wr_cycle[ 1375] = 1'b1;  addr_rom[ 1375]='h00000050;  wr_data_rom[ 1375]='h000003c4;
    rd_cycle[ 1376] = 1'b1;  wr_cycle[ 1376] = 1'b0;  addr_rom[ 1376]='h000007f4;  wr_data_rom[ 1376]='h00000000;
    rd_cycle[ 1377] = 1'b1;  wr_cycle[ 1377] = 1'b0;  addr_rom[ 1377]='h000006f8;  wr_data_rom[ 1377]='h00000000;
    rd_cycle[ 1378] = 1'b1;  wr_cycle[ 1378] = 1'b0;  addr_rom[ 1378]='h000002c0;  wr_data_rom[ 1378]='h00000000;
    rd_cycle[ 1379] = 1'b1;  wr_cycle[ 1379] = 1'b0;  addr_rom[ 1379]='h00000430;  wr_data_rom[ 1379]='h00000000;
    rd_cycle[ 1380] = 1'b1;  wr_cycle[ 1380] = 1'b0;  addr_rom[ 1380]='h00000494;  wr_data_rom[ 1380]='h00000000;
    rd_cycle[ 1381] = 1'b0;  wr_cycle[ 1381] = 1'b1;  addr_rom[ 1381]='h000002d4;  wr_data_rom[ 1381]='h000003d7;
    rd_cycle[ 1382] = 1'b0;  wr_cycle[ 1382] = 1'b1;  addr_rom[ 1382]='h0000014c;  wr_data_rom[ 1382]='h00000048;
    rd_cycle[ 1383] = 1'b1;  wr_cycle[ 1383] = 1'b0;  addr_rom[ 1383]='h000002c8;  wr_data_rom[ 1383]='h00000000;
    rd_cycle[ 1384] = 1'b1;  wr_cycle[ 1384] = 1'b0;  addr_rom[ 1384]='h0000055c;  wr_data_rom[ 1384]='h00000000;
    rd_cycle[ 1385] = 1'b0;  wr_cycle[ 1385] = 1'b1;  addr_rom[ 1385]='h0000024c;  wr_data_rom[ 1385]='h0000030c;
    rd_cycle[ 1386] = 1'b1;  wr_cycle[ 1386] = 1'b0;  addr_rom[ 1386]='h00000600;  wr_data_rom[ 1386]='h00000000;
    rd_cycle[ 1387] = 1'b0;  wr_cycle[ 1387] = 1'b1;  addr_rom[ 1387]='h0000047c;  wr_data_rom[ 1387]='h000000d2;
    rd_cycle[ 1388] = 1'b0;  wr_cycle[ 1388] = 1'b1;  addr_rom[ 1388]='h00000258;  wr_data_rom[ 1388]='h000004df;
    rd_cycle[ 1389] = 1'b1;  wr_cycle[ 1389] = 1'b0;  addr_rom[ 1389]='h00000654;  wr_data_rom[ 1389]='h00000000;
    rd_cycle[ 1390] = 1'b0;  wr_cycle[ 1390] = 1'b1;  addr_rom[ 1390]='h00000780;  wr_data_rom[ 1390]='h00000509;
    rd_cycle[ 1391] = 1'b0;  wr_cycle[ 1391] = 1'b1;  addr_rom[ 1391]='h0000007c;  wr_data_rom[ 1391]='h000002a8;
    rd_cycle[ 1392] = 1'b1;  wr_cycle[ 1392] = 1'b0;  addr_rom[ 1392]='h00000568;  wr_data_rom[ 1392]='h00000000;
    rd_cycle[ 1393] = 1'b0;  wr_cycle[ 1393] = 1'b1;  addr_rom[ 1393]='h00000724;  wr_data_rom[ 1393]='h000000b6;
    rd_cycle[ 1394] = 1'b0;  wr_cycle[ 1394] = 1'b1;  addr_rom[ 1394]='h000002d4;  wr_data_rom[ 1394]='h000002b4;
    rd_cycle[ 1395] = 1'b0;  wr_cycle[ 1395] = 1'b1;  addr_rom[ 1395]='h000006c4;  wr_data_rom[ 1395]='h0000062e;
    rd_cycle[ 1396] = 1'b0;  wr_cycle[ 1396] = 1'b1;  addr_rom[ 1396]='h00000558;  wr_data_rom[ 1396]='h0000017b;
    rd_cycle[ 1397] = 1'b1;  wr_cycle[ 1397] = 1'b0;  addr_rom[ 1397]='h0000067c;  wr_data_rom[ 1397]='h00000000;
    rd_cycle[ 1398] = 1'b1;  wr_cycle[ 1398] = 1'b0;  addr_rom[ 1398]='h000005e0;  wr_data_rom[ 1398]='h00000000;
    rd_cycle[ 1399] = 1'b1;  wr_cycle[ 1399] = 1'b0;  addr_rom[ 1399]='h000002b8;  wr_data_rom[ 1399]='h00000000;
    rd_cycle[ 1400] = 1'b0;  wr_cycle[ 1400] = 1'b1;  addr_rom[ 1400]='h00000148;  wr_data_rom[ 1400]='h00000240;
    rd_cycle[ 1401] = 1'b1;  wr_cycle[ 1401] = 1'b0;  addr_rom[ 1401]='h00000060;  wr_data_rom[ 1401]='h00000000;
    rd_cycle[ 1402] = 1'b1;  wr_cycle[ 1402] = 1'b0;  addr_rom[ 1402]='h000001d4;  wr_data_rom[ 1402]='h00000000;
    rd_cycle[ 1403] = 1'b1;  wr_cycle[ 1403] = 1'b0;  addr_rom[ 1403]='h00000164;  wr_data_rom[ 1403]='h00000000;
    rd_cycle[ 1404] = 1'b0;  wr_cycle[ 1404] = 1'b1;  addr_rom[ 1404]='h0000074c;  wr_data_rom[ 1404]='h00000508;
    rd_cycle[ 1405] = 1'b0;  wr_cycle[ 1405] = 1'b1;  addr_rom[ 1405]='h00000704;  wr_data_rom[ 1405]='h00000424;
    rd_cycle[ 1406] = 1'b1;  wr_cycle[ 1406] = 1'b0;  addr_rom[ 1406]='h000004e4;  wr_data_rom[ 1406]='h00000000;
    rd_cycle[ 1407] = 1'b1;  wr_cycle[ 1407] = 1'b0;  addr_rom[ 1407]='h00000434;  wr_data_rom[ 1407]='h00000000;
    rd_cycle[ 1408] = 1'b0;  wr_cycle[ 1408] = 1'b1;  addr_rom[ 1408]='h000005dc;  wr_data_rom[ 1408]='h0000062c;
    rd_cycle[ 1409] = 1'b1;  wr_cycle[ 1409] = 1'b0;  addr_rom[ 1409]='h00000378;  wr_data_rom[ 1409]='h00000000;
    rd_cycle[ 1410] = 1'b1;  wr_cycle[ 1410] = 1'b0;  addr_rom[ 1410]='h000002c4;  wr_data_rom[ 1410]='h00000000;
    rd_cycle[ 1411] = 1'b0;  wr_cycle[ 1411] = 1'b1;  addr_rom[ 1411]='h00000668;  wr_data_rom[ 1411]='h000002dd;
    rd_cycle[ 1412] = 1'b0;  wr_cycle[ 1412] = 1'b1;  addr_rom[ 1412]='h000005e4;  wr_data_rom[ 1412]='h000006f4;
    rd_cycle[ 1413] = 1'b1;  wr_cycle[ 1413] = 1'b0;  addr_rom[ 1413]='h0000046c;  wr_data_rom[ 1413]='h00000000;
    rd_cycle[ 1414] = 1'b0;  wr_cycle[ 1414] = 1'b1;  addr_rom[ 1414]='h000006ec;  wr_data_rom[ 1414]='h00000396;
    rd_cycle[ 1415] = 1'b1;  wr_cycle[ 1415] = 1'b0;  addr_rom[ 1415]='h00000568;  wr_data_rom[ 1415]='h00000000;
    rd_cycle[ 1416] = 1'b0;  wr_cycle[ 1416] = 1'b1;  addr_rom[ 1416]='h00000284;  wr_data_rom[ 1416]='h000002bd;
    rd_cycle[ 1417] = 1'b1;  wr_cycle[ 1417] = 1'b0;  addr_rom[ 1417]='h00000284;  wr_data_rom[ 1417]='h00000000;
    rd_cycle[ 1418] = 1'b0;  wr_cycle[ 1418] = 1'b1;  addr_rom[ 1418]='h0000061c;  wr_data_rom[ 1418]='h0000009c;
    rd_cycle[ 1419] = 1'b1;  wr_cycle[ 1419] = 1'b0;  addr_rom[ 1419]='h00000440;  wr_data_rom[ 1419]='h00000000;
    rd_cycle[ 1420] = 1'b0;  wr_cycle[ 1420] = 1'b1;  addr_rom[ 1420]='h00000434;  wr_data_rom[ 1420]='h000003aa;
    rd_cycle[ 1421] = 1'b1;  wr_cycle[ 1421] = 1'b0;  addr_rom[ 1421]='h00000488;  wr_data_rom[ 1421]='h00000000;
    rd_cycle[ 1422] = 1'b1;  wr_cycle[ 1422] = 1'b0;  addr_rom[ 1422]='h000003bc;  wr_data_rom[ 1422]='h00000000;
    rd_cycle[ 1423] = 1'b0;  wr_cycle[ 1423] = 1'b1;  addr_rom[ 1423]='h0000061c;  wr_data_rom[ 1423]='h0000027b;
    rd_cycle[ 1424] = 1'b0;  wr_cycle[ 1424] = 1'b1;  addr_rom[ 1424]='h00000528;  wr_data_rom[ 1424]='h000001b8;
    rd_cycle[ 1425] = 1'b1;  wr_cycle[ 1425] = 1'b0;  addr_rom[ 1425]='h000006ac;  wr_data_rom[ 1425]='h00000000;
    rd_cycle[ 1426] = 1'b0;  wr_cycle[ 1426] = 1'b1;  addr_rom[ 1426]='h00000658;  wr_data_rom[ 1426]='h00000149;
    rd_cycle[ 1427] = 1'b1;  wr_cycle[ 1427] = 1'b0;  addr_rom[ 1427]='h000004c0;  wr_data_rom[ 1427]='h00000000;
    rd_cycle[ 1428] = 1'b1;  wr_cycle[ 1428] = 1'b0;  addr_rom[ 1428]='h0000051c;  wr_data_rom[ 1428]='h00000000;
    rd_cycle[ 1429] = 1'b0;  wr_cycle[ 1429] = 1'b1;  addr_rom[ 1429]='h000002d0;  wr_data_rom[ 1429]='h0000067b;
    rd_cycle[ 1430] = 1'b1;  wr_cycle[ 1430] = 1'b0;  addr_rom[ 1430]='h000000c0;  wr_data_rom[ 1430]='h00000000;
    rd_cycle[ 1431] = 1'b1;  wr_cycle[ 1431] = 1'b0;  addr_rom[ 1431]='h000004bc;  wr_data_rom[ 1431]='h00000000;
    rd_cycle[ 1432] = 1'b0;  wr_cycle[ 1432] = 1'b1;  addr_rom[ 1432]='h00000510;  wr_data_rom[ 1432]='h000006f1;
    rd_cycle[ 1433] = 1'b0;  wr_cycle[ 1433] = 1'b1;  addr_rom[ 1433]='h000006b4;  wr_data_rom[ 1433]='h0000018a;
    rd_cycle[ 1434] = 1'b0;  wr_cycle[ 1434] = 1'b1;  addr_rom[ 1434]='h000000f0;  wr_data_rom[ 1434]='h000000be;
    rd_cycle[ 1435] = 1'b0;  wr_cycle[ 1435] = 1'b1;  addr_rom[ 1435]='h00000334;  wr_data_rom[ 1435]='h000004fe;
    rd_cycle[ 1436] = 1'b0;  wr_cycle[ 1436] = 1'b1;  addr_rom[ 1436]='h00000540;  wr_data_rom[ 1436]='h0000063a;
    rd_cycle[ 1437] = 1'b1;  wr_cycle[ 1437] = 1'b0;  addr_rom[ 1437]='h000005fc;  wr_data_rom[ 1437]='h00000000;
    rd_cycle[ 1438] = 1'b1;  wr_cycle[ 1438] = 1'b0;  addr_rom[ 1438]='h00000770;  wr_data_rom[ 1438]='h00000000;
    rd_cycle[ 1439] = 1'b1;  wr_cycle[ 1439] = 1'b0;  addr_rom[ 1439]='h000002a8;  wr_data_rom[ 1439]='h00000000;
    rd_cycle[ 1440] = 1'b1;  wr_cycle[ 1440] = 1'b0;  addr_rom[ 1440]='h000007e0;  wr_data_rom[ 1440]='h00000000;
    rd_cycle[ 1441] = 1'b1;  wr_cycle[ 1441] = 1'b0;  addr_rom[ 1441]='h00000130;  wr_data_rom[ 1441]='h00000000;
    rd_cycle[ 1442] = 1'b0;  wr_cycle[ 1442] = 1'b1;  addr_rom[ 1442]='h00000550;  wr_data_rom[ 1442]='h00000304;
    rd_cycle[ 1443] = 1'b0;  wr_cycle[ 1443] = 1'b1;  addr_rom[ 1443]='h00000460;  wr_data_rom[ 1443]='h00000691;
    rd_cycle[ 1444] = 1'b0;  wr_cycle[ 1444] = 1'b1;  addr_rom[ 1444]='h00000168;  wr_data_rom[ 1444]='h000004cf;
    rd_cycle[ 1445] = 1'b0;  wr_cycle[ 1445] = 1'b1;  addr_rom[ 1445]='h00000790;  wr_data_rom[ 1445]='h000002f5;
    rd_cycle[ 1446] = 1'b1;  wr_cycle[ 1446] = 1'b0;  addr_rom[ 1446]='h00000638;  wr_data_rom[ 1446]='h00000000;
    rd_cycle[ 1447] = 1'b0;  wr_cycle[ 1447] = 1'b1;  addr_rom[ 1447]='h00000550;  wr_data_rom[ 1447]='h000005a1;
    rd_cycle[ 1448] = 1'b0;  wr_cycle[ 1448] = 1'b1;  addr_rom[ 1448]='h00000144;  wr_data_rom[ 1448]='h000004a6;
    rd_cycle[ 1449] = 1'b0;  wr_cycle[ 1449] = 1'b1;  addr_rom[ 1449]='h000001a0;  wr_data_rom[ 1449]='h0000029d;
    rd_cycle[ 1450] = 1'b1;  wr_cycle[ 1450] = 1'b0;  addr_rom[ 1450]='h00000270;  wr_data_rom[ 1450]='h00000000;
    rd_cycle[ 1451] = 1'b1;  wr_cycle[ 1451] = 1'b0;  addr_rom[ 1451]='h00000598;  wr_data_rom[ 1451]='h00000000;
    rd_cycle[ 1452] = 1'b1;  wr_cycle[ 1452] = 1'b0;  addr_rom[ 1452]='h0000066c;  wr_data_rom[ 1452]='h00000000;
    rd_cycle[ 1453] = 1'b0;  wr_cycle[ 1453] = 1'b1;  addr_rom[ 1453]='h000001dc;  wr_data_rom[ 1453]='h00000170;
    rd_cycle[ 1454] = 1'b1;  wr_cycle[ 1454] = 1'b0;  addr_rom[ 1454]='h00000724;  wr_data_rom[ 1454]='h00000000;
    rd_cycle[ 1455] = 1'b0;  wr_cycle[ 1455] = 1'b1;  addr_rom[ 1455]='h00000430;  wr_data_rom[ 1455]='h0000066f;
    rd_cycle[ 1456] = 1'b1;  wr_cycle[ 1456] = 1'b0;  addr_rom[ 1456]='h000006a0;  wr_data_rom[ 1456]='h00000000;
    rd_cycle[ 1457] = 1'b1;  wr_cycle[ 1457] = 1'b0;  addr_rom[ 1457]='h00000468;  wr_data_rom[ 1457]='h00000000;
    rd_cycle[ 1458] = 1'b1;  wr_cycle[ 1458] = 1'b0;  addr_rom[ 1458]='h00000544;  wr_data_rom[ 1458]='h00000000;
    rd_cycle[ 1459] = 1'b0;  wr_cycle[ 1459] = 1'b1;  addr_rom[ 1459]='h000004d0;  wr_data_rom[ 1459]='h0000020c;
    rd_cycle[ 1460] = 1'b1;  wr_cycle[ 1460] = 1'b0;  addr_rom[ 1460]='h000006dc;  wr_data_rom[ 1460]='h00000000;
    rd_cycle[ 1461] = 1'b1;  wr_cycle[ 1461] = 1'b0;  addr_rom[ 1461]='h00000758;  wr_data_rom[ 1461]='h00000000;
    rd_cycle[ 1462] = 1'b1;  wr_cycle[ 1462] = 1'b0;  addr_rom[ 1462]='h00000108;  wr_data_rom[ 1462]='h00000000;
    rd_cycle[ 1463] = 1'b1;  wr_cycle[ 1463] = 1'b0;  addr_rom[ 1463]='h00000014;  wr_data_rom[ 1463]='h00000000;
    rd_cycle[ 1464] = 1'b1;  wr_cycle[ 1464] = 1'b0;  addr_rom[ 1464]='h000007dc;  wr_data_rom[ 1464]='h00000000;
    rd_cycle[ 1465] = 1'b1;  wr_cycle[ 1465] = 1'b0;  addr_rom[ 1465]='h0000008c;  wr_data_rom[ 1465]='h00000000;
    rd_cycle[ 1466] = 1'b1;  wr_cycle[ 1466] = 1'b0;  addr_rom[ 1466]='h000002b0;  wr_data_rom[ 1466]='h00000000;
    rd_cycle[ 1467] = 1'b0;  wr_cycle[ 1467] = 1'b1;  addr_rom[ 1467]='h0000007c;  wr_data_rom[ 1467]='h0000006d;
    rd_cycle[ 1468] = 1'b1;  wr_cycle[ 1468] = 1'b0;  addr_rom[ 1468]='h00000338;  wr_data_rom[ 1468]='h00000000;
    rd_cycle[ 1469] = 1'b1;  wr_cycle[ 1469] = 1'b0;  addr_rom[ 1469]='h00000020;  wr_data_rom[ 1469]='h00000000;
    rd_cycle[ 1470] = 1'b1;  wr_cycle[ 1470] = 1'b0;  addr_rom[ 1470]='h00000114;  wr_data_rom[ 1470]='h00000000;
    rd_cycle[ 1471] = 1'b0;  wr_cycle[ 1471] = 1'b1;  addr_rom[ 1471]='h0000069c;  wr_data_rom[ 1471]='h00000664;
    rd_cycle[ 1472] = 1'b0;  wr_cycle[ 1472] = 1'b1;  addr_rom[ 1472]='h00000158;  wr_data_rom[ 1472]='h000000e2;
    rd_cycle[ 1473] = 1'b0;  wr_cycle[ 1473] = 1'b1;  addr_rom[ 1473]='h000005c4;  wr_data_rom[ 1473]='h000002a9;
    rd_cycle[ 1474] = 1'b1;  wr_cycle[ 1474] = 1'b0;  addr_rom[ 1474]='h00000390;  wr_data_rom[ 1474]='h00000000;
    rd_cycle[ 1475] = 1'b1;  wr_cycle[ 1475] = 1'b0;  addr_rom[ 1475]='h000006f4;  wr_data_rom[ 1475]='h00000000;
    rd_cycle[ 1476] = 1'b1;  wr_cycle[ 1476] = 1'b0;  addr_rom[ 1476]='h000003a0;  wr_data_rom[ 1476]='h00000000;
    rd_cycle[ 1477] = 1'b1;  wr_cycle[ 1477] = 1'b0;  addr_rom[ 1477]='h00000638;  wr_data_rom[ 1477]='h00000000;
    rd_cycle[ 1478] = 1'b1;  wr_cycle[ 1478] = 1'b0;  addr_rom[ 1478]='h000002c0;  wr_data_rom[ 1478]='h00000000;
    rd_cycle[ 1479] = 1'b0;  wr_cycle[ 1479] = 1'b1;  addr_rom[ 1479]='h00000548;  wr_data_rom[ 1479]='h00000106;
    rd_cycle[ 1480] = 1'b0;  wr_cycle[ 1480] = 1'b1;  addr_rom[ 1480]='h000004d0;  wr_data_rom[ 1480]='h000000bb;
    rd_cycle[ 1481] = 1'b0;  wr_cycle[ 1481] = 1'b1;  addr_rom[ 1481]='h0000066c;  wr_data_rom[ 1481]='h000003a3;
    rd_cycle[ 1482] = 1'b1;  wr_cycle[ 1482] = 1'b0;  addr_rom[ 1482]='h00000448;  wr_data_rom[ 1482]='h00000000;
    rd_cycle[ 1483] = 1'b1;  wr_cycle[ 1483] = 1'b0;  addr_rom[ 1483]='h00000678;  wr_data_rom[ 1483]='h00000000;
    rd_cycle[ 1484] = 1'b1;  wr_cycle[ 1484] = 1'b0;  addr_rom[ 1484]='h00000780;  wr_data_rom[ 1484]='h00000000;
    rd_cycle[ 1485] = 1'b1;  wr_cycle[ 1485] = 1'b0;  addr_rom[ 1485]='h00000624;  wr_data_rom[ 1485]='h00000000;
    rd_cycle[ 1486] = 1'b1;  wr_cycle[ 1486] = 1'b0;  addr_rom[ 1486]='h000005fc;  wr_data_rom[ 1486]='h00000000;
    rd_cycle[ 1487] = 1'b0;  wr_cycle[ 1487] = 1'b1;  addr_rom[ 1487]='h00000758;  wr_data_rom[ 1487]='h00000387;
    rd_cycle[ 1488] = 1'b0;  wr_cycle[ 1488] = 1'b1;  addr_rom[ 1488]='h0000036c;  wr_data_rom[ 1488]='h0000051a;
    rd_cycle[ 1489] = 1'b1;  wr_cycle[ 1489] = 1'b0;  addr_rom[ 1489]='h00000318;  wr_data_rom[ 1489]='h00000000;
    rd_cycle[ 1490] = 1'b0;  wr_cycle[ 1490] = 1'b1;  addr_rom[ 1490]='h0000054c;  wr_data_rom[ 1490]='h00000559;
    rd_cycle[ 1491] = 1'b1;  wr_cycle[ 1491] = 1'b0;  addr_rom[ 1491]='h00000704;  wr_data_rom[ 1491]='h00000000;
    rd_cycle[ 1492] = 1'b0;  wr_cycle[ 1492] = 1'b1;  addr_rom[ 1492]='h000005c4;  wr_data_rom[ 1492]='h00000540;
    rd_cycle[ 1493] = 1'b0;  wr_cycle[ 1493] = 1'b1;  addr_rom[ 1493]='h0000011c;  wr_data_rom[ 1493]='h000006b1;
    rd_cycle[ 1494] = 1'b1;  wr_cycle[ 1494] = 1'b0;  addr_rom[ 1494]='h000001c4;  wr_data_rom[ 1494]='h00000000;
    rd_cycle[ 1495] = 1'b0;  wr_cycle[ 1495] = 1'b1;  addr_rom[ 1495]='h00000560;  wr_data_rom[ 1495]='h00000735;
    rd_cycle[ 1496] = 1'b0;  wr_cycle[ 1496] = 1'b1;  addr_rom[ 1496]='h00000200;  wr_data_rom[ 1496]='h000006de;
    rd_cycle[ 1497] = 1'b0;  wr_cycle[ 1497] = 1'b1;  addr_rom[ 1497]='h00000610;  wr_data_rom[ 1497]='h000002d5;
    rd_cycle[ 1498] = 1'b1;  wr_cycle[ 1498] = 1'b0;  addr_rom[ 1498]='h000001d0;  wr_data_rom[ 1498]='h00000000;
    rd_cycle[ 1499] = 1'b1;  wr_cycle[ 1499] = 1'b0;  addr_rom[ 1499]='h000000d8;  wr_data_rom[ 1499]='h00000000;
    rd_cycle[ 1500] = 1'b1;  wr_cycle[ 1500] = 1'b0;  addr_rom[ 1500]='h000004e0;  wr_data_rom[ 1500]='h00000000;
    rd_cycle[ 1501] = 1'b1;  wr_cycle[ 1501] = 1'b0;  addr_rom[ 1501]='h00000608;  wr_data_rom[ 1501]='h00000000;
    rd_cycle[ 1502] = 1'b1;  wr_cycle[ 1502] = 1'b0;  addr_rom[ 1502]='h000007ac;  wr_data_rom[ 1502]='h00000000;
    rd_cycle[ 1503] = 1'b0;  wr_cycle[ 1503] = 1'b1;  addr_rom[ 1503]='h0000020c;  wr_data_rom[ 1503]='h00000549;
    rd_cycle[ 1504] = 1'b1;  wr_cycle[ 1504] = 1'b0;  addr_rom[ 1504]='h00000634;  wr_data_rom[ 1504]='h00000000;
    rd_cycle[ 1505] = 1'b0;  wr_cycle[ 1505] = 1'b1;  addr_rom[ 1505]='h00000458;  wr_data_rom[ 1505]='h0000075b;
    rd_cycle[ 1506] = 1'b0;  wr_cycle[ 1506] = 1'b1;  addr_rom[ 1506]='h00000570;  wr_data_rom[ 1506]='h000001d3;
    rd_cycle[ 1507] = 1'b1;  wr_cycle[ 1507] = 1'b0;  addr_rom[ 1507]='h000004dc;  wr_data_rom[ 1507]='h00000000;
    rd_cycle[ 1508] = 1'b1;  wr_cycle[ 1508] = 1'b0;  addr_rom[ 1508]='h000004cc;  wr_data_rom[ 1508]='h00000000;
    rd_cycle[ 1509] = 1'b0;  wr_cycle[ 1509] = 1'b1;  addr_rom[ 1509]='h000002c0;  wr_data_rom[ 1509]='h000000a9;
    rd_cycle[ 1510] = 1'b1;  wr_cycle[ 1510] = 1'b0;  addr_rom[ 1510]='h000003c0;  wr_data_rom[ 1510]='h00000000;
    rd_cycle[ 1511] = 1'b0;  wr_cycle[ 1511] = 1'b1;  addr_rom[ 1511]='h00000048;  wr_data_rom[ 1511]='h00000345;
    rd_cycle[ 1512] = 1'b0;  wr_cycle[ 1512] = 1'b1;  addr_rom[ 1512]='h00000710;  wr_data_rom[ 1512]='h0000079c;
    rd_cycle[ 1513] = 1'b0;  wr_cycle[ 1513] = 1'b1;  addr_rom[ 1513]='h000005f0;  wr_data_rom[ 1513]='h000005c2;
    rd_cycle[ 1514] = 1'b0;  wr_cycle[ 1514] = 1'b1;  addr_rom[ 1514]='h000001c0;  wr_data_rom[ 1514]='h00000071;
    rd_cycle[ 1515] = 1'b1;  wr_cycle[ 1515] = 1'b0;  addr_rom[ 1515]='h000001a0;  wr_data_rom[ 1515]='h00000000;
    rd_cycle[ 1516] = 1'b1;  wr_cycle[ 1516] = 1'b0;  addr_rom[ 1516]='h000005cc;  wr_data_rom[ 1516]='h00000000;
    rd_cycle[ 1517] = 1'b0;  wr_cycle[ 1517] = 1'b1;  addr_rom[ 1517]='h00000190;  wr_data_rom[ 1517]='h0000008e;
    rd_cycle[ 1518] = 1'b1;  wr_cycle[ 1518] = 1'b0;  addr_rom[ 1518]='h00000508;  wr_data_rom[ 1518]='h00000000;
    rd_cycle[ 1519] = 1'b0;  wr_cycle[ 1519] = 1'b1;  addr_rom[ 1519]='h000002ac;  wr_data_rom[ 1519]='h0000035f;
    rd_cycle[ 1520] = 1'b1;  wr_cycle[ 1520] = 1'b0;  addr_rom[ 1520]='h00000670;  wr_data_rom[ 1520]='h00000000;
    rd_cycle[ 1521] = 1'b0;  wr_cycle[ 1521] = 1'b1;  addr_rom[ 1521]='h00000334;  wr_data_rom[ 1521]='h00000709;
    rd_cycle[ 1522] = 1'b1;  wr_cycle[ 1522] = 1'b0;  addr_rom[ 1522]='h00000650;  wr_data_rom[ 1522]='h00000000;
    rd_cycle[ 1523] = 1'b0;  wr_cycle[ 1523] = 1'b1;  addr_rom[ 1523]='h00000678;  wr_data_rom[ 1523]='h00000000;
    rd_cycle[ 1524] = 1'b1;  wr_cycle[ 1524] = 1'b0;  addr_rom[ 1524]='h00000680;  wr_data_rom[ 1524]='h00000000;
    rd_cycle[ 1525] = 1'b0;  wr_cycle[ 1525] = 1'b1;  addr_rom[ 1525]='h000001fc;  wr_data_rom[ 1525]='h000004c5;
    rd_cycle[ 1526] = 1'b1;  wr_cycle[ 1526] = 1'b0;  addr_rom[ 1526]='h000007a4;  wr_data_rom[ 1526]='h00000000;
    rd_cycle[ 1527] = 1'b0;  wr_cycle[ 1527] = 1'b1;  addr_rom[ 1527]='h000005c4;  wr_data_rom[ 1527]='h000004cc;
    rd_cycle[ 1528] = 1'b0;  wr_cycle[ 1528] = 1'b1;  addr_rom[ 1528]='h000006c8;  wr_data_rom[ 1528]='h00000003;
    rd_cycle[ 1529] = 1'b1;  wr_cycle[ 1529] = 1'b0;  addr_rom[ 1529]='h00000040;  wr_data_rom[ 1529]='h00000000;
    rd_cycle[ 1530] = 1'b0;  wr_cycle[ 1530] = 1'b1;  addr_rom[ 1530]='h00000584;  wr_data_rom[ 1530]='h00000547;
    rd_cycle[ 1531] = 1'b0;  wr_cycle[ 1531] = 1'b1;  addr_rom[ 1531]='h0000028c;  wr_data_rom[ 1531]='h00000595;
    rd_cycle[ 1532] = 1'b1;  wr_cycle[ 1532] = 1'b0;  addr_rom[ 1532]='h00000754;  wr_data_rom[ 1532]='h00000000;
    rd_cycle[ 1533] = 1'b1;  wr_cycle[ 1533] = 1'b0;  addr_rom[ 1533]='h00000650;  wr_data_rom[ 1533]='h00000000;
    rd_cycle[ 1534] = 1'b0;  wr_cycle[ 1534] = 1'b1;  addr_rom[ 1534]='h00000334;  wr_data_rom[ 1534]='h000005a6;
    rd_cycle[ 1535] = 1'b1;  wr_cycle[ 1535] = 1'b0;  addr_rom[ 1535]='h00000258;  wr_data_rom[ 1535]='h00000000;
    rd_cycle[ 1536] = 1'b0;  wr_cycle[ 1536] = 1'b1;  addr_rom[ 1536]='h000004ec;  wr_data_rom[ 1536]='h00000403;
    rd_cycle[ 1537] = 1'b1;  wr_cycle[ 1537] = 1'b0;  addr_rom[ 1537]='h00000008;  wr_data_rom[ 1537]='h00000000;
    rd_cycle[ 1538] = 1'b1;  wr_cycle[ 1538] = 1'b0;  addr_rom[ 1538]='h00000178;  wr_data_rom[ 1538]='h00000000;
    rd_cycle[ 1539] = 1'b0;  wr_cycle[ 1539] = 1'b1;  addr_rom[ 1539]='h00000628;  wr_data_rom[ 1539]='h000005c1;
    rd_cycle[ 1540] = 1'b0;  wr_cycle[ 1540] = 1'b1;  addr_rom[ 1540]='h0000040c;  wr_data_rom[ 1540]='h000001db;
    rd_cycle[ 1541] = 1'b1;  wr_cycle[ 1541] = 1'b0;  addr_rom[ 1541]='h000000f4;  wr_data_rom[ 1541]='h00000000;
    rd_cycle[ 1542] = 1'b1;  wr_cycle[ 1542] = 1'b0;  addr_rom[ 1542]='h00000568;  wr_data_rom[ 1542]='h00000000;
    rd_cycle[ 1543] = 1'b1;  wr_cycle[ 1543] = 1'b0;  addr_rom[ 1543]='h000005c8;  wr_data_rom[ 1543]='h00000000;
    rd_cycle[ 1544] = 1'b0;  wr_cycle[ 1544] = 1'b1;  addr_rom[ 1544]='h00000334;  wr_data_rom[ 1544]='h00000528;
    rd_cycle[ 1545] = 1'b1;  wr_cycle[ 1545] = 1'b0;  addr_rom[ 1545]='h00000410;  wr_data_rom[ 1545]='h00000000;
    rd_cycle[ 1546] = 1'b0;  wr_cycle[ 1546] = 1'b1;  addr_rom[ 1546]='h00000010;  wr_data_rom[ 1546]='h000007ca;
    rd_cycle[ 1547] = 1'b1;  wr_cycle[ 1547] = 1'b0;  addr_rom[ 1547]='h00000468;  wr_data_rom[ 1547]='h00000000;
    rd_cycle[ 1548] = 1'b1;  wr_cycle[ 1548] = 1'b0;  addr_rom[ 1548]='h000002d4;  wr_data_rom[ 1548]='h00000000;
    rd_cycle[ 1549] = 1'b1;  wr_cycle[ 1549] = 1'b0;  addr_rom[ 1549]='h00000608;  wr_data_rom[ 1549]='h00000000;
    rd_cycle[ 1550] = 1'b1;  wr_cycle[ 1550] = 1'b0;  addr_rom[ 1550]='h00000240;  wr_data_rom[ 1550]='h00000000;
    rd_cycle[ 1551] = 1'b0;  wr_cycle[ 1551] = 1'b1;  addr_rom[ 1551]='h00000668;  wr_data_rom[ 1551]='h0000033f;
    rd_cycle[ 1552] = 1'b0;  wr_cycle[ 1552] = 1'b1;  addr_rom[ 1552]='h00000250;  wr_data_rom[ 1552]='h0000056f;
    rd_cycle[ 1553] = 1'b0;  wr_cycle[ 1553] = 1'b1;  addr_rom[ 1553]='h00000220;  wr_data_rom[ 1553]='h0000018c;
    rd_cycle[ 1554] = 1'b0;  wr_cycle[ 1554] = 1'b1;  addr_rom[ 1554]='h0000047c;  wr_data_rom[ 1554]='h00000628;
    rd_cycle[ 1555] = 1'b1;  wr_cycle[ 1555] = 1'b0;  addr_rom[ 1555]='h00000250;  wr_data_rom[ 1555]='h00000000;
    rd_cycle[ 1556] = 1'b1;  wr_cycle[ 1556] = 1'b0;  addr_rom[ 1556]='h00000794;  wr_data_rom[ 1556]='h00000000;
    rd_cycle[ 1557] = 1'b0;  wr_cycle[ 1557] = 1'b1;  addr_rom[ 1557]='h00000608;  wr_data_rom[ 1557]='h0000021c;
    rd_cycle[ 1558] = 1'b0;  wr_cycle[ 1558] = 1'b1;  addr_rom[ 1558]='h000004a0;  wr_data_rom[ 1558]='h0000065d;
    rd_cycle[ 1559] = 1'b1;  wr_cycle[ 1559] = 1'b0;  addr_rom[ 1559]='h000005cc;  wr_data_rom[ 1559]='h00000000;
    rd_cycle[ 1560] = 1'b1;  wr_cycle[ 1560] = 1'b0;  addr_rom[ 1560]='h00000604;  wr_data_rom[ 1560]='h00000000;
    rd_cycle[ 1561] = 1'b1;  wr_cycle[ 1561] = 1'b0;  addr_rom[ 1561]='h000001ac;  wr_data_rom[ 1561]='h00000000;
    rd_cycle[ 1562] = 1'b1;  wr_cycle[ 1562] = 1'b0;  addr_rom[ 1562]='h0000047c;  wr_data_rom[ 1562]='h00000000;
    rd_cycle[ 1563] = 1'b0;  wr_cycle[ 1563] = 1'b1;  addr_rom[ 1563]='h00000034;  wr_data_rom[ 1563]='h000006e5;
    rd_cycle[ 1564] = 1'b0;  wr_cycle[ 1564] = 1'b1;  addr_rom[ 1564]='h000006a4;  wr_data_rom[ 1564]='h00000689;
    rd_cycle[ 1565] = 1'b1;  wr_cycle[ 1565] = 1'b0;  addr_rom[ 1565]='h000007d4;  wr_data_rom[ 1565]='h00000000;
    rd_cycle[ 1566] = 1'b0;  wr_cycle[ 1566] = 1'b1;  addr_rom[ 1566]='h000000dc;  wr_data_rom[ 1566]='h000002af;
    rd_cycle[ 1567] = 1'b0;  wr_cycle[ 1567] = 1'b1;  addr_rom[ 1567]='h00000090;  wr_data_rom[ 1567]='h0000068a;
    rd_cycle[ 1568] = 1'b0;  wr_cycle[ 1568] = 1'b1;  addr_rom[ 1568]='h00000610;  wr_data_rom[ 1568]='h00000665;
    rd_cycle[ 1569] = 1'b0;  wr_cycle[ 1569] = 1'b1;  addr_rom[ 1569]='h00000648;  wr_data_rom[ 1569]='h00000574;
    rd_cycle[ 1570] = 1'b1;  wr_cycle[ 1570] = 1'b0;  addr_rom[ 1570]='h000007b4;  wr_data_rom[ 1570]='h00000000;
    rd_cycle[ 1571] = 1'b1;  wr_cycle[ 1571] = 1'b0;  addr_rom[ 1571]='h00000474;  wr_data_rom[ 1571]='h00000000;
    rd_cycle[ 1572] = 1'b0;  wr_cycle[ 1572] = 1'b1;  addr_rom[ 1572]='h000003e8;  wr_data_rom[ 1572]='h0000033c;
    rd_cycle[ 1573] = 1'b0;  wr_cycle[ 1573] = 1'b1;  addr_rom[ 1573]='h00000270;  wr_data_rom[ 1573]='h0000068c;
    rd_cycle[ 1574] = 1'b1;  wr_cycle[ 1574] = 1'b0;  addr_rom[ 1574]='h000004fc;  wr_data_rom[ 1574]='h00000000;
    rd_cycle[ 1575] = 1'b1;  wr_cycle[ 1575] = 1'b0;  addr_rom[ 1575]='h0000069c;  wr_data_rom[ 1575]='h00000000;
    rd_cycle[ 1576] = 1'b1;  wr_cycle[ 1576] = 1'b0;  addr_rom[ 1576]='h00000294;  wr_data_rom[ 1576]='h00000000;
    rd_cycle[ 1577] = 1'b0;  wr_cycle[ 1577] = 1'b1;  addr_rom[ 1577]='h00000184;  wr_data_rom[ 1577]='h00000390;
    rd_cycle[ 1578] = 1'b1;  wr_cycle[ 1578] = 1'b0;  addr_rom[ 1578]='h000007ec;  wr_data_rom[ 1578]='h00000000;
    rd_cycle[ 1579] = 1'b1;  wr_cycle[ 1579] = 1'b0;  addr_rom[ 1579]='h00000480;  wr_data_rom[ 1579]='h00000000;
    rd_cycle[ 1580] = 1'b0;  wr_cycle[ 1580] = 1'b1;  addr_rom[ 1580]='h00000280;  wr_data_rom[ 1580]='h00000402;
    rd_cycle[ 1581] = 1'b0;  wr_cycle[ 1581] = 1'b1;  addr_rom[ 1581]='h00000578;  wr_data_rom[ 1581]='h00000098;
    rd_cycle[ 1582] = 1'b0;  wr_cycle[ 1582] = 1'b1;  addr_rom[ 1582]='h00000110;  wr_data_rom[ 1582]='h0000013b;
    rd_cycle[ 1583] = 1'b0;  wr_cycle[ 1583] = 1'b1;  addr_rom[ 1583]='h000002a8;  wr_data_rom[ 1583]='h0000011c;
    rd_cycle[ 1584] = 1'b0;  wr_cycle[ 1584] = 1'b1;  addr_rom[ 1584]='h00000200;  wr_data_rom[ 1584]='h000002c9;
    rd_cycle[ 1585] = 1'b1;  wr_cycle[ 1585] = 1'b0;  addr_rom[ 1585]='h000006e0;  wr_data_rom[ 1585]='h00000000;
    rd_cycle[ 1586] = 1'b0;  wr_cycle[ 1586] = 1'b1;  addr_rom[ 1586]='h0000023c;  wr_data_rom[ 1586]='h0000043d;
    rd_cycle[ 1587] = 1'b0;  wr_cycle[ 1587] = 1'b1;  addr_rom[ 1587]='h000003c0;  wr_data_rom[ 1587]='h0000042a;
    rd_cycle[ 1588] = 1'b0;  wr_cycle[ 1588] = 1'b1;  addr_rom[ 1588]='h00000320;  wr_data_rom[ 1588]='h000002d9;
    rd_cycle[ 1589] = 1'b0;  wr_cycle[ 1589] = 1'b1;  addr_rom[ 1589]='h000004f0;  wr_data_rom[ 1589]='h00000302;
    rd_cycle[ 1590] = 1'b1;  wr_cycle[ 1590] = 1'b0;  addr_rom[ 1590]='h000001a8;  wr_data_rom[ 1590]='h00000000;
    rd_cycle[ 1591] = 1'b1;  wr_cycle[ 1591] = 1'b0;  addr_rom[ 1591]='h000000fc;  wr_data_rom[ 1591]='h00000000;
    rd_cycle[ 1592] = 1'b0;  wr_cycle[ 1592] = 1'b1;  addr_rom[ 1592]='h0000073c;  wr_data_rom[ 1592]='h00000523;
    rd_cycle[ 1593] = 1'b1;  wr_cycle[ 1593] = 1'b0;  addr_rom[ 1593]='h000003d0;  wr_data_rom[ 1593]='h00000000;
    rd_cycle[ 1594] = 1'b1;  wr_cycle[ 1594] = 1'b0;  addr_rom[ 1594]='h00000024;  wr_data_rom[ 1594]='h00000000;
    rd_cycle[ 1595] = 1'b0;  wr_cycle[ 1595] = 1'b1;  addr_rom[ 1595]='h00000510;  wr_data_rom[ 1595]='h0000059a;
    rd_cycle[ 1596] = 1'b0;  wr_cycle[ 1596] = 1'b1;  addr_rom[ 1596]='h00000074;  wr_data_rom[ 1596]='h00000753;
    rd_cycle[ 1597] = 1'b1;  wr_cycle[ 1597] = 1'b0;  addr_rom[ 1597]='h00000610;  wr_data_rom[ 1597]='h00000000;
    rd_cycle[ 1598] = 1'b1;  wr_cycle[ 1598] = 1'b0;  addr_rom[ 1598]='h000007cc;  wr_data_rom[ 1598]='h00000000;
    rd_cycle[ 1599] = 1'b1;  wr_cycle[ 1599] = 1'b0;  addr_rom[ 1599]='h00000388;  wr_data_rom[ 1599]='h00000000;
    rd_cycle[ 1600] = 1'b0;  wr_cycle[ 1600] = 1'b1;  addr_rom[ 1600]='h000006d0;  wr_data_rom[ 1600]='h000004b7;
    rd_cycle[ 1601] = 1'b0;  wr_cycle[ 1601] = 1'b1;  addr_rom[ 1601]='h00000540;  wr_data_rom[ 1601]='h0000020c;
    rd_cycle[ 1602] = 1'b1;  wr_cycle[ 1602] = 1'b0;  addr_rom[ 1602]='h00000678;  wr_data_rom[ 1602]='h00000000;
    rd_cycle[ 1603] = 1'b0;  wr_cycle[ 1603] = 1'b1;  addr_rom[ 1603]='h000002ec;  wr_data_rom[ 1603]='h0000025d;
    rd_cycle[ 1604] = 1'b0;  wr_cycle[ 1604] = 1'b1;  addr_rom[ 1604]='h00000468;  wr_data_rom[ 1604]='h000004f4;
    rd_cycle[ 1605] = 1'b0;  wr_cycle[ 1605] = 1'b1;  addr_rom[ 1605]='h00000004;  wr_data_rom[ 1605]='h0000065b;
    rd_cycle[ 1606] = 1'b1;  wr_cycle[ 1606] = 1'b0;  addr_rom[ 1606]='h000001d0;  wr_data_rom[ 1606]='h00000000;
    rd_cycle[ 1607] = 1'b0;  wr_cycle[ 1607] = 1'b1;  addr_rom[ 1607]='h00000088;  wr_data_rom[ 1607]='h0000062f;
    rd_cycle[ 1608] = 1'b1;  wr_cycle[ 1608] = 1'b0;  addr_rom[ 1608]='h000004a0;  wr_data_rom[ 1608]='h00000000;
    rd_cycle[ 1609] = 1'b1;  wr_cycle[ 1609] = 1'b0;  addr_rom[ 1609]='h0000017c;  wr_data_rom[ 1609]='h00000000;
    rd_cycle[ 1610] = 1'b1;  wr_cycle[ 1610] = 1'b0;  addr_rom[ 1610]='h000005d4;  wr_data_rom[ 1610]='h00000000;
    rd_cycle[ 1611] = 1'b0;  wr_cycle[ 1611] = 1'b1;  addr_rom[ 1611]='h00000468;  wr_data_rom[ 1611]='h00000112;
    rd_cycle[ 1612] = 1'b0;  wr_cycle[ 1612] = 1'b1;  addr_rom[ 1612]='h000007dc;  wr_data_rom[ 1612]='h00000379;
    rd_cycle[ 1613] = 1'b0;  wr_cycle[ 1613] = 1'b1;  addr_rom[ 1613]='h00000114;  wr_data_rom[ 1613]='h000002ef;
    rd_cycle[ 1614] = 1'b1;  wr_cycle[ 1614] = 1'b0;  addr_rom[ 1614]='h00000178;  wr_data_rom[ 1614]='h00000000;
    rd_cycle[ 1615] = 1'b1;  wr_cycle[ 1615] = 1'b0;  addr_rom[ 1615]='h00000384;  wr_data_rom[ 1615]='h00000000;
    rd_cycle[ 1616] = 1'b1;  wr_cycle[ 1616] = 1'b0;  addr_rom[ 1616]='h00000338;  wr_data_rom[ 1616]='h00000000;
    rd_cycle[ 1617] = 1'b1;  wr_cycle[ 1617] = 1'b0;  addr_rom[ 1617]='h000000dc;  wr_data_rom[ 1617]='h00000000;
    rd_cycle[ 1618] = 1'b0;  wr_cycle[ 1618] = 1'b1;  addr_rom[ 1618]='h00000068;  wr_data_rom[ 1618]='h00000399;
    rd_cycle[ 1619] = 1'b0;  wr_cycle[ 1619] = 1'b1;  addr_rom[ 1619]='h000004bc;  wr_data_rom[ 1619]='h00000591;
    rd_cycle[ 1620] = 1'b0;  wr_cycle[ 1620] = 1'b1;  addr_rom[ 1620]='h000001d0;  wr_data_rom[ 1620]='h000000a0;
    rd_cycle[ 1621] = 1'b1;  wr_cycle[ 1621] = 1'b0;  addr_rom[ 1621]='h000001b0;  wr_data_rom[ 1621]='h00000000;
    rd_cycle[ 1622] = 1'b1;  wr_cycle[ 1622] = 1'b0;  addr_rom[ 1622]='h000006ac;  wr_data_rom[ 1622]='h00000000;
    rd_cycle[ 1623] = 1'b0;  wr_cycle[ 1623] = 1'b1;  addr_rom[ 1623]='h00000400;  wr_data_rom[ 1623]='h00000382;
    rd_cycle[ 1624] = 1'b0;  wr_cycle[ 1624] = 1'b1;  addr_rom[ 1624]='h00000138;  wr_data_rom[ 1624]='h0000061a;
    rd_cycle[ 1625] = 1'b1;  wr_cycle[ 1625] = 1'b0;  addr_rom[ 1625]='h0000001c;  wr_data_rom[ 1625]='h00000000;
    rd_cycle[ 1626] = 1'b0;  wr_cycle[ 1626] = 1'b1;  addr_rom[ 1626]='h000001b8;  wr_data_rom[ 1626]='h000004c5;
    rd_cycle[ 1627] = 1'b0;  wr_cycle[ 1627] = 1'b1;  addr_rom[ 1627]='h00000360;  wr_data_rom[ 1627]='h000005dd;
    rd_cycle[ 1628] = 1'b1;  wr_cycle[ 1628] = 1'b0;  addr_rom[ 1628]='h00000554;  wr_data_rom[ 1628]='h00000000;
    rd_cycle[ 1629] = 1'b0;  wr_cycle[ 1629] = 1'b1;  addr_rom[ 1629]='h000007c0;  wr_data_rom[ 1629]='h00000690;
    rd_cycle[ 1630] = 1'b0;  wr_cycle[ 1630] = 1'b1;  addr_rom[ 1630]='h000005f4;  wr_data_rom[ 1630]='h0000053f;
    rd_cycle[ 1631] = 1'b1;  wr_cycle[ 1631] = 1'b0;  addr_rom[ 1631]='h00000030;  wr_data_rom[ 1631]='h00000000;
    rd_cycle[ 1632] = 1'b1;  wr_cycle[ 1632] = 1'b0;  addr_rom[ 1632]='h00000074;  wr_data_rom[ 1632]='h00000000;
    rd_cycle[ 1633] = 1'b0;  wr_cycle[ 1633] = 1'b1;  addr_rom[ 1633]='h000000ec;  wr_data_rom[ 1633]='h000004c0;
    rd_cycle[ 1634] = 1'b0;  wr_cycle[ 1634] = 1'b1;  addr_rom[ 1634]='h00000394;  wr_data_rom[ 1634]='h00000555;
    rd_cycle[ 1635] = 1'b1;  wr_cycle[ 1635] = 1'b0;  addr_rom[ 1635]='h00000098;  wr_data_rom[ 1635]='h00000000;
    rd_cycle[ 1636] = 1'b0;  wr_cycle[ 1636] = 1'b1;  addr_rom[ 1636]='h00000078;  wr_data_rom[ 1636]='h00000058;
    rd_cycle[ 1637] = 1'b1;  wr_cycle[ 1637] = 1'b0;  addr_rom[ 1637]='h00000550;  wr_data_rom[ 1637]='h00000000;
    rd_cycle[ 1638] = 1'b0;  wr_cycle[ 1638] = 1'b1;  addr_rom[ 1638]='h000000ec;  wr_data_rom[ 1638]='h000003d7;
    rd_cycle[ 1639] = 1'b0;  wr_cycle[ 1639] = 1'b1;  addr_rom[ 1639]='h00000628;  wr_data_rom[ 1639]='h00000005;
    rd_cycle[ 1640] = 1'b0;  wr_cycle[ 1640] = 1'b1;  addr_rom[ 1640]='h00000194;  wr_data_rom[ 1640]='h00000012;
    rd_cycle[ 1641] = 1'b1;  wr_cycle[ 1641] = 1'b0;  addr_rom[ 1641]='h000005b8;  wr_data_rom[ 1641]='h00000000;
    rd_cycle[ 1642] = 1'b0;  wr_cycle[ 1642] = 1'b1;  addr_rom[ 1642]='h00000128;  wr_data_rom[ 1642]='h0000011a;
    rd_cycle[ 1643] = 1'b1;  wr_cycle[ 1643] = 1'b0;  addr_rom[ 1643]='h00000450;  wr_data_rom[ 1643]='h00000000;
    rd_cycle[ 1644] = 1'b0;  wr_cycle[ 1644] = 1'b1;  addr_rom[ 1644]='h00000414;  wr_data_rom[ 1644]='h000001c2;
    rd_cycle[ 1645] = 1'b1;  wr_cycle[ 1645] = 1'b0;  addr_rom[ 1645]='h00000048;  wr_data_rom[ 1645]='h00000000;
    rd_cycle[ 1646] = 1'b0;  wr_cycle[ 1646] = 1'b1;  addr_rom[ 1646]='h000007b8;  wr_data_rom[ 1646]='h00000362;
    rd_cycle[ 1647] = 1'b0;  wr_cycle[ 1647] = 1'b1;  addr_rom[ 1647]='h00000728;  wr_data_rom[ 1647]='h0000054e;
    rd_cycle[ 1648] = 1'b1;  wr_cycle[ 1648] = 1'b0;  addr_rom[ 1648]='h00000270;  wr_data_rom[ 1648]='h00000000;
    rd_cycle[ 1649] = 1'b1;  wr_cycle[ 1649] = 1'b0;  addr_rom[ 1649]='h00000538;  wr_data_rom[ 1649]='h00000000;
    rd_cycle[ 1650] = 1'b0;  wr_cycle[ 1650] = 1'b1;  addr_rom[ 1650]='h000000f8;  wr_data_rom[ 1650]='h000007e9;
    rd_cycle[ 1651] = 1'b0;  wr_cycle[ 1651] = 1'b1;  addr_rom[ 1651]='h00000708;  wr_data_rom[ 1651]='h00000184;
    rd_cycle[ 1652] = 1'b1;  wr_cycle[ 1652] = 1'b0;  addr_rom[ 1652]='h00000634;  wr_data_rom[ 1652]='h00000000;
    rd_cycle[ 1653] = 1'b0;  wr_cycle[ 1653] = 1'b1;  addr_rom[ 1653]='h0000055c;  wr_data_rom[ 1653]='h00000750;
    rd_cycle[ 1654] = 1'b0;  wr_cycle[ 1654] = 1'b1;  addr_rom[ 1654]='h000003c8;  wr_data_rom[ 1654]='h000003d3;
    rd_cycle[ 1655] = 1'b1;  wr_cycle[ 1655] = 1'b0;  addr_rom[ 1655]='h00000234;  wr_data_rom[ 1655]='h00000000;
    rd_cycle[ 1656] = 1'b0;  wr_cycle[ 1656] = 1'b1;  addr_rom[ 1656]='h0000042c;  wr_data_rom[ 1656]='h000003f7;
    rd_cycle[ 1657] = 1'b0;  wr_cycle[ 1657] = 1'b1;  addr_rom[ 1657]='h000007cc;  wr_data_rom[ 1657]='h000007fd;
    rd_cycle[ 1658] = 1'b1;  wr_cycle[ 1658] = 1'b0;  addr_rom[ 1658]='h00000650;  wr_data_rom[ 1658]='h00000000;
    rd_cycle[ 1659] = 1'b1;  wr_cycle[ 1659] = 1'b0;  addr_rom[ 1659]='h00000360;  wr_data_rom[ 1659]='h00000000;
    rd_cycle[ 1660] = 1'b1;  wr_cycle[ 1660] = 1'b0;  addr_rom[ 1660]='h000002bc;  wr_data_rom[ 1660]='h00000000;
    rd_cycle[ 1661] = 1'b0;  wr_cycle[ 1661] = 1'b1;  addr_rom[ 1661]='h0000007c;  wr_data_rom[ 1661]='h00000526;
    rd_cycle[ 1662] = 1'b0;  wr_cycle[ 1662] = 1'b1;  addr_rom[ 1662]='h00000068;  wr_data_rom[ 1662]='h00000765;
    rd_cycle[ 1663] = 1'b0;  wr_cycle[ 1663] = 1'b1;  addr_rom[ 1663]='h000002bc;  wr_data_rom[ 1663]='h000002b4;
    rd_cycle[ 1664] = 1'b1;  wr_cycle[ 1664] = 1'b0;  addr_rom[ 1664]='h00000180;  wr_data_rom[ 1664]='h00000000;
    rd_cycle[ 1665] = 1'b1;  wr_cycle[ 1665] = 1'b0;  addr_rom[ 1665]='h00000418;  wr_data_rom[ 1665]='h00000000;
    rd_cycle[ 1666] = 1'b1;  wr_cycle[ 1666] = 1'b0;  addr_rom[ 1666]='h000007a0;  wr_data_rom[ 1666]='h00000000;
    rd_cycle[ 1667] = 1'b1;  wr_cycle[ 1667] = 1'b0;  addr_rom[ 1667]='h000006f8;  wr_data_rom[ 1667]='h00000000;
    rd_cycle[ 1668] = 1'b1;  wr_cycle[ 1668] = 1'b0;  addr_rom[ 1668]='h00000768;  wr_data_rom[ 1668]='h00000000;
    rd_cycle[ 1669] = 1'b0;  wr_cycle[ 1669] = 1'b1;  addr_rom[ 1669]='h00000660;  wr_data_rom[ 1669]='h0000031d;
    rd_cycle[ 1670] = 1'b1;  wr_cycle[ 1670] = 1'b0;  addr_rom[ 1670]='h0000028c;  wr_data_rom[ 1670]='h00000000;
    rd_cycle[ 1671] = 1'b0;  wr_cycle[ 1671] = 1'b1;  addr_rom[ 1671]='h00000044;  wr_data_rom[ 1671]='h00000266;
    rd_cycle[ 1672] = 1'b1;  wr_cycle[ 1672] = 1'b0;  addr_rom[ 1672]='h0000028c;  wr_data_rom[ 1672]='h00000000;
    rd_cycle[ 1673] = 1'b0;  wr_cycle[ 1673] = 1'b1;  addr_rom[ 1673]='h0000013c;  wr_data_rom[ 1673]='h0000005d;
    rd_cycle[ 1674] = 1'b1;  wr_cycle[ 1674] = 1'b0;  addr_rom[ 1674]='h000000e8;  wr_data_rom[ 1674]='h00000000;
    rd_cycle[ 1675] = 1'b1;  wr_cycle[ 1675] = 1'b0;  addr_rom[ 1675]='h0000075c;  wr_data_rom[ 1675]='h00000000;
    rd_cycle[ 1676] = 1'b0;  wr_cycle[ 1676] = 1'b1;  addr_rom[ 1676]='h000000c4;  wr_data_rom[ 1676]='h000000b5;
    rd_cycle[ 1677] = 1'b1;  wr_cycle[ 1677] = 1'b0;  addr_rom[ 1677]='h00000150;  wr_data_rom[ 1677]='h00000000;
    rd_cycle[ 1678] = 1'b0;  wr_cycle[ 1678] = 1'b1;  addr_rom[ 1678]='h00000788;  wr_data_rom[ 1678]='h00000234;
    rd_cycle[ 1679] = 1'b1;  wr_cycle[ 1679] = 1'b0;  addr_rom[ 1679]='h0000039c;  wr_data_rom[ 1679]='h00000000;
    rd_cycle[ 1680] = 1'b1;  wr_cycle[ 1680] = 1'b0;  addr_rom[ 1680]='h000003dc;  wr_data_rom[ 1680]='h00000000;
    rd_cycle[ 1681] = 1'b0;  wr_cycle[ 1681] = 1'b1;  addr_rom[ 1681]='h0000012c;  wr_data_rom[ 1681]='h0000033b;
    rd_cycle[ 1682] = 1'b1;  wr_cycle[ 1682] = 1'b0;  addr_rom[ 1682]='h00000614;  wr_data_rom[ 1682]='h00000000;
    rd_cycle[ 1683] = 1'b0;  wr_cycle[ 1683] = 1'b1;  addr_rom[ 1683]='h00000134;  wr_data_rom[ 1683]='h00000639;
    rd_cycle[ 1684] = 1'b1;  wr_cycle[ 1684] = 1'b0;  addr_rom[ 1684]='h000000cc;  wr_data_rom[ 1684]='h00000000;
    rd_cycle[ 1685] = 1'b1;  wr_cycle[ 1685] = 1'b0;  addr_rom[ 1685]='h000003cc;  wr_data_rom[ 1685]='h00000000;
    rd_cycle[ 1686] = 1'b1;  wr_cycle[ 1686] = 1'b0;  addr_rom[ 1686]='h000000c0;  wr_data_rom[ 1686]='h00000000;
    rd_cycle[ 1687] = 1'b0;  wr_cycle[ 1687] = 1'b1;  addr_rom[ 1687]='h00000648;  wr_data_rom[ 1687]='h0000072b;
    rd_cycle[ 1688] = 1'b0;  wr_cycle[ 1688] = 1'b1;  addr_rom[ 1688]='h000007ac;  wr_data_rom[ 1688]='h000003e9;
    rd_cycle[ 1689] = 1'b1;  wr_cycle[ 1689] = 1'b0;  addr_rom[ 1689]='h000004f4;  wr_data_rom[ 1689]='h00000000;
    rd_cycle[ 1690] = 1'b0;  wr_cycle[ 1690] = 1'b1;  addr_rom[ 1690]='h00000468;  wr_data_rom[ 1690]='h0000028b;
    rd_cycle[ 1691] = 1'b1;  wr_cycle[ 1691] = 1'b0;  addr_rom[ 1691]='h000003a0;  wr_data_rom[ 1691]='h00000000;
    rd_cycle[ 1692] = 1'b1;  wr_cycle[ 1692] = 1'b0;  addr_rom[ 1692]='h000000e4;  wr_data_rom[ 1692]='h00000000;
    rd_cycle[ 1693] = 1'b0;  wr_cycle[ 1693] = 1'b1;  addr_rom[ 1693]='h00000510;  wr_data_rom[ 1693]='h000002f7;
    rd_cycle[ 1694] = 1'b1;  wr_cycle[ 1694] = 1'b0;  addr_rom[ 1694]='h00000768;  wr_data_rom[ 1694]='h00000000;
    rd_cycle[ 1695] = 1'b1;  wr_cycle[ 1695] = 1'b0;  addr_rom[ 1695]='h000005a8;  wr_data_rom[ 1695]='h00000000;
    rd_cycle[ 1696] = 1'b0;  wr_cycle[ 1696] = 1'b1;  addr_rom[ 1696]='h0000024c;  wr_data_rom[ 1696]='h00000203;
    rd_cycle[ 1697] = 1'b0;  wr_cycle[ 1697] = 1'b1;  addr_rom[ 1697]='h0000077c;  wr_data_rom[ 1697]='h00000022;
    rd_cycle[ 1698] = 1'b0;  wr_cycle[ 1698] = 1'b1;  addr_rom[ 1698]='h00000270;  wr_data_rom[ 1698]='h000001f9;
    rd_cycle[ 1699] = 1'b1;  wr_cycle[ 1699] = 1'b0;  addr_rom[ 1699]='h0000027c;  wr_data_rom[ 1699]='h00000000;
    rd_cycle[ 1700] = 1'b1;  wr_cycle[ 1700] = 1'b0;  addr_rom[ 1700]='h00000740;  wr_data_rom[ 1700]='h00000000;
    rd_cycle[ 1701] = 1'b0;  wr_cycle[ 1701] = 1'b1;  addr_rom[ 1701]='h00000668;  wr_data_rom[ 1701]='h000002ae;
    rd_cycle[ 1702] = 1'b0;  wr_cycle[ 1702] = 1'b1;  addr_rom[ 1702]='h00000230;  wr_data_rom[ 1702]='h0000019e;
    rd_cycle[ 1703] = 1'b0;  wr_cycle[ 1703] = 1'b1;  addr_rom[ 1703]='h00000710;  wr_data_rom[ 1703]='h0000022c;
    rd_cycle[ 1704] = 1'b1;  wr_cycle[ 1704] = 1'b0;  addr_rom[ 1704]='h0000030c;  wr_data_rom[ 1704]='h00000000;
    rd_cycle[ 1705] = 1'b1;  wr_cycle[ 1705] = 1'b0;  addr_rom[ 1705]='h00000194;  wr_data_rom[ 1705]='h00000000;
    rd_cycle[ 1706] = 1'b1;  wr_cycle[ 1706] = 1'b0;  addr_rom[ 1706]='h00000438;  wr_data_rom[ 1706]='h00000000;
    rd_cycle[ 1707] = 1'b1;  wr_cycle[ 1707] = 1'b0;  addr_rom[ 1707]='h000001d0;  wr_data_rom[ 1707]='h00000000;
    rd_cycle[ 1708] = 1'b1;  wr_cycle[ 1708] = 1'b0;  addr_rom[ 1708]='h00000478;  wr_data_rom[ 1708]='h00000000;
    rd_cycle[ 1709] = 1'b1;  wr_cycle[ 1709] = 1'b0;  addr_rom[ 1709]='h00000130;  wr_data_rom[ 1709]='h00000000;
    rd_cycle[ 1710] = 1'b1;  wr_cycle[ 1710] = 1'b0;  addr_rom[ 1710]='h00000324;  wr_data_rom[ 1710]='h00000000;
    rd_cycle[ 1711] = 1'b1;  wr_cycle[ 1711] = 1'b0;  addr_rom[ 1711]='h00000284;  wr_data_rom[ 1711]='h00000000;
    rd_cycle[ 1712] = 1'b1;  wr_cycle[ 1712] = 1'b0;  addr_rom[ 1712]='h000003c0;  wr_data_rom[ 1712]='h00000000;
    rd_cycle[ 1713] = 1'b0;  wr_cycle[ 1713] = 1'b1;  addr_rom[ 1713]='h0000014c;  wr_data_rom[ 1713]='h00000273;
    rd_cycle[ 1714] = 1'b1;  wr_cycle[ 1714] = 1'b0;  addr_rom[ 1714]='h000007b8;  wr_data_rom[ 1714]='h00000000;
    rd_cycle[ 1715] = 1'b1;  wr_cycle[ 1715] = 1'b0;  addr_rom[ 1715]='h000007a4;  wr_data_rom[ 1715]='h00000000;
    rd_cycle[ 1716] = 1'b0;  wr_cycle[ 1716] = 1'b1;  addr_rom[ 1716]='h000006c0;  wr_data_rom[ 1716]='h00000487;
    rd_cycle[ 1717] = 1'b1;  wr_cycle[ 1717] = 1'b0;  addr_rom[ 1717]='h00000740;  wr_data_rom[ 1717]='h00000000;
    rd_cycle[ 1718] = 1'b1;  wr_cycle[ 1718] = 1'b0;  addr_rom[ 1718]='h000003b0;  wr_data_rom[ 1718]='h00000000;
    rd_cycle[ 1719] = 1'b1;  wr_cycle[ 1719] = 1'b0;  addr_rom[ 1719]='h0000016c;  wr_data_rom[ 1719]='h00000000;
    rd_cycle[ 1720] = 1'b0;  wr_cycle[ 1720] = 1'b1;  addr_rom[ 1720]='h00000448;  wr_data_rom[ 1720]='h00000791;
    rd_cycle[ 1721] = 1'b1;  wr_cycle[ 1721] = 1'b0;  addr_rom[ 1721]='h00000548;  wr_data_rom[ 1721]='h00000000;
    rd_cycle[ 1722] = 1'b1;  wr_cycle[ 1722] = 1'b0;  addr_rom[ 1722]='h00000670;  wr_data_rom[ 1722]='h00000000;
    rd_cycle[ 1723] = 1'b1;  wr_cycle[ 1723] = 1'b0;  addr_rom[ 1723]='h0000059c;  wr_data_rom[ 1723]='h00000000;
    rd_cycle[ 1724] = 1'b1;  wr_cycle[ 1724] = 1'b0;  addr_rom[ 1724]='h00000010;  wr_data_rom[ 1724]='h00000000;
    rd_cycle[ 1725] = 1'b1;  wr_cycle[ 1725] = 1'b0;  addr_rom[ 1725]='h00000454;  wr_data_rom[ 1725]='h00000000;
    rd_cycle[ 1726] = 1'b1;  wr_cycle[ 1726] = 1'b0;  addr_rom[ 1726]='h000007f4;  wr_data_rom[ 1726]='h00000000;
    rd_cycle[ 1727] = 1'b1;  wr_cycle[ 1727] = 1'b0;  addr_rom[ 1727]='h0000050c;  wr_data_rom[ 1727]='h00000000;
    rd_cycle[ 1728] = 1'b0;  wr_cycle[ 1728] = 1'b1;  addr_rom[ 1728]='h000006e0;  wr_data_rom[ 1728]='h00000693;
    rd_cycle[ 1729] = 1'b1;  wr_cycle[ 1729] = 1'b0;  addr_rom[ 1729]='h000001f4;  wr_data_rom[ 1729]='h00000000;
    rd_cycle[ 1730] = 1'b1;  wr_cycle[ 1730] = 1'b0;  addr_rom[ 1730]='h000001e4;  wr_data_rom[ 1730]='h00000000;
    rd_cycle[ 1731] = 1'b0;  wr_cycle[ 1731] = 1'b1;  addr_rom[ 1731]='h00000148;  wr_data_rom[ 1731]='h000001cb;
    rd_cycle[ 1732] = 1'b1;  wr_cycle[ 1732] = 1'b0;  addr_rom[ 1732]='h000003c8;  wr_data_rom[ 1732]='h00000000;
    rd_cycle[ 1733] = 1'b1;  wr_cycle[ 1733] = 1'b0;  addr_rom[ 1733]='h00000240;  wr_data_rom[ 1733]='h00000000;
    rd_cycle[ 1734] = 1'b1;  wr_cycle[ 1734] = 1'b0;  addr_rom[ 1734]='h00000090;  wr_data_rom[ 1734]='h00000000;
    rd_cycle[ 1735] = 1'b1;  wr_cycle[ 1735] = 1'b0;  addr_rom[ 1735]='h000007e8;  wr_data_rom[ 1735]='h00000000;
    rd_cycle[ 1736] = 1'b0;  wr_cycle[ 1736] = 1'b1;  addr_rom[ 1736]='h00000018;  wr_data_rom[ 1736]='h0000027c;
    rd_cycle[ 1737] = 1'b1;  wr_cycle[ 1737] = 1'b0;  addr_rom[ 1737]='h000003fc;  wr_data_rom[ 1737]='h00000000;
    rd_cycle[ 1738] = 1'b0;  wr_cycle[ 1738] = 1'b1;  addr_rom[ 1738]='h00000738;  wr_data_rom[ 1738]='h0000052e;
    rd_cycle[ 1739] = 1'b1;  wr_cycle[ 1739] = 1'b0;  addr_rom[ 1739]='h00000774;  wr_data_rom[ 1739]='h00000000;
    rd_cycle[ 1740] = 1'b0;  wr_cycle[ 1740] = 1'b1;  addr_rom[ 1740]='h000004a8;  wr_data_rom[ 1740]='h0000071b;
    rd_cycle[ 1741] = 1'b1;  wr_cycle[ 1741] = 1'b0;  addr_rom[ 1741]='h000006dc;  wr_data_rom[ 1741]='h00000000;
    rd_cycle[ 1742] = 1'b1;  wr_cycle[ 1742] = 1'b0;  addr_rom[ 1742]='h000003f4;  wr_data_rom[ 1742]='h00000000;
    rd_cycle[ 1743] = 1'b1;  wr_cycle[ 1743] = 1'b0;  addr_rom[ 1743]='h0000055c;  wr_data_rom[ 1743]='h00000000;
    rd_cycle[ 1744] = 1'b0;  wr_cycle[ 1744] = 1'b1;  addr_rom[ 1744]='h000002c4;  wr_data_rom[ 1744]='h000004f8;
    rd_cycle[ 1745] = 1'b1;  wr_cycle[ 1745] = 1'b0;  addr_rom[ 1745]='h00000788;  wr_data_rom[ 1745]='h00000000;
    rd_cycle[ 1746] = 1'b1;  wr_cycle[ 1746] = 1'b0;  addr_rom[ 1746]='h00000730;  wr_data_rom[ 1746]='h00000000;
    rd_cycle[ 1747] = 1'b1;  wr_cycle[ 1747] = 1'b0;  addr_rom[ 1747]='h00000594;  wr_data_rom[ 1747]='h00000000;
    rd_cycle[ 1748] = 1'b1;  wr_cycle[ 1748] = 1'b0;  addr_rom[ 1748]='h000001b0;  wr_data_rom[ 1748]='h00000000;
    rd_cycle[ 1749] = 1'b0;  wr_cycle[ 1749] = 1'b1;  addr_rom[ 1749]='h0000015c;  wr_data_rom[ 1749]='h00000089;
    rd_cycle[ 1750] = 1'b0;  wr_cycle[ 1750] = 1'b1;  addr_rom[ 1750]='h00000170;  wr_data_rom[ 1750]='h000005d1;
    rd_cycle[ 1751] = 1'b1;  wr_cycle[ 1751] = 1'b0;  addr_rom[ 1751]='h00000220;  wr_data_rom[ 1751]='h00000000;
    rd_cycle[ 1752] = 1'b1;  wr_cycle[ 1752] = 1'b0;  addr_rom[ 1752]='h000001f8;  wr_data_rom[ 1752]='h00000000;
    rd_cycle[ 1753] = 1'b1;  wr_cycle[ 1753] = 1'b0;  addr_rom[ 1753]='h000000a8;  wr_data_rom[ 1753]='h00000000;
    rd_cycle[ 1754] = 1'b0;  wr_cycle[ 1754] = 1'b1;  addr_rom[ 1754]='h000003f8;  wr_data_rom[ 1754]='h00000243;
    rd_cycle[ 1755] = 1'b0;  wr_cycle[ 1755] = 1'b1;  addr_rom[ 1755]='h00000374;  wr_data_rom[ 1755]='h0000067a;
    rd_cycle[ 1756] = 1'b0;  wr_cycle[ 1756] = 1'b1;  addr_rom[ 1756]='h00000004;  wr_data_rom[ 1756]='h000001e6;
    rd_cycle[ 1757] = 1'b0;  wr_cycle[ 1757] = 1'b1;  addr_rom[ 1757]='h000005d4;  wr_data_rom[ 1757]='h00000553;
    rd_cycle[ 1758] = 1'b0;  wr_cycle[ 1758] = 1'b1;  addr_rom[ 1758]='h00000258;  wr_data_rom[ 1758]='h000002b2;
    rd_cycle[ 1759] = 1'b1;  wr_cycle[ 1759] = 1'b0;  addr_rom[ 1759]='h0000046c;  wr_data_rom[ 1759]='h00000000;
    rd_cycle[ 1760] = 1'b1;  wr_cycle[ 1760] = 1'b0;  addr_rom[ 1760]='h00000250;  wr_data_rom[ 1760]='h00000000;
    rd_cycle[ 1761] = 1'b0;  wr_cycle[ 1761] = 1'b1;  addr_rom[ 1761]='h00000228;  wr_data_rom[ 1761]='h00000432;
    rd_cycle[ 1762] = 1'b1;  wr_cycle[ 1762] = 1'b0;  addr_rom[ 1762]='h00000414;  wr_data_rom[ 1762]='h00000000;
    rd_cycle[ 1763] = 1'b0;  wr_cycle[ 1763] = 1'b1;  addr_rom[ 1763]='h000002c8;  wr_data_rom[ 1763]='h000002f7;
    rd_cycle[ 1764] = 1'b1;  wr_cycle[ 1764] = 1'b0;  addr_rom[ 1764]='h00000784;  wr_data_rom[ 1764]='h00000000;
    rd_cycle[ 1765] = 1'b0;  wr_cycle[ 1765] = 1'b1;  addr_rom[ 1765]='h000001c4;  wr_data_rom[ 1765]='h000005fd;
    rd_cycle[ 1766] = 1'b0;  wr_cycle[ 1766] = 1'b1;  addr_rom[ 1766]='h000001e8;  wr_data_rom[ 1766]='h00000514;
    rd_cycle[ 1767] = 1'b0;  wr_cycle[ 1767] = 1'b1;  addr_rom[ 1767]='h00000328;  wr_data_rom[ 1767]='h0000059d;
    rd_cycle[ 1768] = 1'b0;  wr_cycle[ 1768] = 1'b1;  addr_rom[ 1768]='h0000009c;  wr_data_rom[ 1768]='h00000533;
    rd_cycle[ 1769] = 1'b0;  wr_cycle[ 1769] = 1'b1;  addr_rom[ 1769]='h00000188;  wr_data_rom[ 1769]='h0000065e;
    rd_cycle[ 1770] = 1'b0;  wr_cycle[ 1770] = 1'b1;  addr_rom[ 1770]='h00000318;  wr_data_rom[ 1770]='h000003fa;
    rd_cycle[ 1771] = 1'b0;  wr_cycle[ 1771] = 1'b1;  addr_rom[ 1771]='h00000624;  wr_data_rom[ 1771]='h000004fc;
    rd_cycle[ 1772] = 1'b1;  wr_cycle[ 1772] = 1'b0;  addr_rom[ 1772]='h000002f8;  wr_data_rom[ 1772]='h00000000;
    rd_cycle[ 1773] = 1'b0;  wr_cycle[ 1773] = 1'b1;  addr_rom[ 1773]='h000004f0;  wr_data_rom[ 1773]='h00000132;
    rd_cycle[ 1774] = 1'b1;  wr_cycle[ 1774] = 1'b0;  addr_rom[ 1774]='h00000250;  wr_data_rom[ 1774]='h00000000;
    rd_cycle[ 1775] = 1'b1;  wr_cycle[ 1775] = 1'b0;  addr_rom[ 1775]='h00000488;  wr_data_rom[ 1775]='h00000000;
    rd_cycle[ 1776] = 1'b0;  wr_cycle[ 1776] = 1'b1;  addr_rom[ 1776]='h00000204;  wr_data_rom[ 1776]='h000002c1;
    rd_cycle[ 1777] = 1'b1;  wr_cycle[ 1777] = 1'b0;  addr_rom[ 1777]='h0000007c;  wr_data_rom[ 1777]='h00000000;
    rd_cycle[ 1778] = 1'b0;  wr_cycle[ 1778] = 1'b1;  addr_rom[ 1778]='h00000060;  wr_data_rom[ 1778]='h00000224;
    rd_cycle[ 1779] = 1'b1;  wr_cycle[ 1779] = 1'b0;  addr_rom[ 1779]='h00000700;  wr_data_rom[ 1779]='h00000000;
    rd_cycle[ 1780] = 1'b0;  wr_cycle[ 1780] = 1'b1;  addr_rom[ 1780]='h00000700;  wr_data_rom[ 1780]='h00000581;
    rd_cycle[ 1781] = 1'b1;  wr_cycle[ 1781] = 1'b0;  addr_rom[ 1781]='h0000021c;  wr_data_rom[ 1781]='h00000000;
    rd_cycle[ 1782] = 1'b0;  wr_cycle[ 1782] = 1'b1;  addr_rom[ 1782]='h0000077c;  wr_data_rom[ 1782]='h000003aa;
    rd_cycle[ 1783] = 1'b1;  wr_cycle[ 1783] = 1'b0;  addr_rom[ 1783]='h000000d8;  wr_data_rom[ 1783]='h00000000;
    rd_cycle[ 1784] = 1'b1;  wr_cycle[ 1784] = 1'b0;  addr_rom[ 1784]='h0000017c;  wr_data_rom[ 1784]='h00000000;
    rd_cycle[ 1785] = 1'b0;  wr_cycle[ 1785] = 1'b1;  addr_rom[ 1785]='h00000034;  wr_data_rom[ 1785]='h00000780;
    rd_cycle[ 1786] = 1'b1;  wr_cycle[ 1786] = 1'b0;  addr_rom[ 1786]='h00000128;  wr_data_rom[ 1786]='h00000000;
    rd_cycle[ 1787] = 1'b0;  wr_cycle[ 1787] = 1'b1;  addr_rom[ 1787]='h000006f0;  wr_data_rom[ 1787]='h00000589;
    rd_cycle[ 1788] = 1'b0;  wr_cycle[ 1788] = 1'b1;  addr_rom[ 1788]='h000003cc;  wr_data_rom[ 1788]='h0000072e;
    rd_cycle[ 1789] = 1'b0;  wr_cycle[ 1789] = 1'b1;  addr_rom[ 1789]='h0000062c;  wr_data_rom[ 1789]='h000003e1;
    rd_cycle[ 1790] = 1'b1;  wr_cycle[ 1790] = 1'b0;  addr_rom[ 1790]='h000002fc;  wr_data_rom[ 1790]='h00000000;
    rd_cycle[ 1791] = 1'b1;  wr_cycle[ 1791] = 1'b0;  addr_rom[ 1791]='h000004f4;  wr_data_rom[ 1791]='h00000000;
    rd_cycle[ 1792] = 1'b0;  wr_cycle[ 1792] = 1'b1;  addr_rom[ 1792]='h00000590;  wr_data_rom[ 1792]='h00000542;
    rd_cycle[ 1793] = 1'b1;  wr_cycle[ 1793] = 1'b0;  addr_rom[ 1793]='h0000014c;  wr_data_rom[ 1793]='h00000000;
    rd_cycle[ 1794] = 1'b0;  wr_cycle[ 1794] = 1'b1;  addr_rom[ 1794]='h0000005c;  wr_data_rom[ 1794]='h000001e2;
    rd_cycle[ 1795] = 1'b1;  wr_cycle[ 1795] = 1'b0;  addr_rom[ 1795]='h0000012c;  wr_data_rom[ 1795]='h00000000;
    rd_cycle[ 1796] = 1'b1;  wr_cycle[ 1796] = 1'b0;  addr_rom[ 1796]='h00000428;  wr_data_rom[ 1796]='h00000000;
    rd_cycle[ 1797] = 1'b1;  wr_cycle[ 1797] = 1'b0;  addr_rom[ 1797]='h000002d4;  wr_data_rom[ 1797]='h00000000;
    rd_cycle[ 1798] = 1'b1;  wr_cycle[ 1798] = 1'b0;  addr_rom[ 1798]='h000000e0;  wr_data_rom[ 1798]='h00000000;
    rd_cycle[ 1799] = 1'b0;  wr_cycle[ 1799] = 1'b1;  addr_rom[ 1799]='h000004e0;  wr_data_rom[ 1799]='h00000484;
    rd_cycle[ 1800] = 1'b1;  wr_cycle[ 1800] = 1'b0;  addr_rom[ 1800]='h0000055c;  wr_data_rom[ 1800]='h00000000;
    rd_cycle[ 1801] = 1'b0;  wr_cycle[ 1801] = 1'b1;  addr_rom[ 1801]='h000006e0;  wr_data_rom[ 1801]='h000002a7;
    rd_cycle[ 1802] = 1'b1;  wr_cycle[ 1802] = 1'b0;  addr_rom[ 1802]='h000000ac;  wr_data_rom[ 1802]='h00000000;
    rd_cycle[ 1803] = 1'b1;  wr_cycle[ 1803] = 1'b0;  addr_rom[ 1803]='h00000538;  wr_data_rom[ 1803]='h00000000;
    rd_cycle[ 1804] = 1'b1;  wr_cycle[ 1804] = 1'b0;  addr_rom[ 1804]='h00000474;  wr_data_rom[ 1804]='h00000000;
    rd_cycle[ 1805] = 1'b0;  wr_cycle[ 1805] = 1'b1;  addr_rom[ 1805]='h0000070c;  wr_data_rom[ 1805]='h0000038e;
    rd_cycle[ 1806] = 1'b0;  wr_cycle[ 1806] = 1'b1;  addr_rom[ 1806]='h0000044c;  wr_data_rom[ 1806]='h00000379;
    rd_cycle[ 1807] = 1'b0;  wr_cycle[ 1807] = 1'b1;  addr_rom[ 1807]='h00000134;  wr_data_rom[ 1807]='h0000011d;
    rd_cycle[ 1808] = 1'b0;  wr_cycle[ 1808] = 1'b1;  addr_rom[ 1808]='h000005c4;  wr_data_rom[ 1808]='h0000071d;
    rd_cycle[ 1809] = 1'b0;  wr_cycle[ 1809] = 1'b1;  addr_rom[ 1809]='h00000780;  wr_data_rom[ 1809]='h00000348;
    rd_cycle[ 1810] = 1'b1;  wr_cycle[ 1810] = 1'b0;  addr_rom[ 1810]='h0000067c;  wr_data_rom[ 1810]='h00000000;
    rd_cycle[ 1811] = 1'b1;  wr_cycle[ 1811] = 1'b0;  addr_rom[ 1811]='h000003a8;  wr_data_rom[ 1811]='h00000000;
    rd_cycle[ 1812] = 1'b0;  wr_cycle[ 1812] = 1'b1;  addr_rom[ 1812]='h00000730;  wr_data_rom[ 1812]='h000000d7;
    rd_cycle[ 1813] = 1'b1;  wr_cycle[ 1813] = 1'b0;  addr_rom[ 1813]='h000007d8;  wr_data_rom[ 1813]='h00000000;
    rd_cycle[ 1814] = 1'b0;  wr_cycle[ 1814] = 1'b1;  addr_rom[ 1814]='h00000180;  wr_data_rom[ 1814]='h0000074e;
    rd_cycle[ 1815] = 1'b0;  wr_cycle[ 1815] = 1'b1;  addr_rom[ 1815]='h000002f8;  wr_data_rom[ 1815]='h0000078b;
    rd_cycle[ 1816] = 1'b1;  wr_cycle[ 1816] = 1'b0;  addr_rom[ 1816]='h00000258;  wr_data_rom[ 1816]='h00000000;
    rd_cycle[ 1817] = 1'b0;  wr_cycle[ 1817] = 1'b1;  addr_rom[ 1817]='h000002fc;  wr_data_rom[ 1817]='h00000215;
    rd_cycle[ 1818] = 1'b1;  wr_cycle[ 1818] = 1'b0;  addr_rom[ 1818]='h00000254;  wr_data_rom[ 1818]='h00000000;
    rd_cycle[ 1819] = 1'b1;  wr_cycle[ 1819] = 1'b0;  addr_rom[ 1819]='h0000054c;  wr_data_rom[ 1819]='h00000000;
    rd_cycle[ 1820] = 1'b1;  wr_cycle[ 1820] = 1'b0;  addr_rom[ 1820]='h000004f0;  wr_data_rom[ 1820]='h00000000;
    rd_cycle[ 1821] = 1'b1;  wr_cycle[ 1821] = 1'b0;  addr_rom[ 1821]='h000006a4;  wr_data_rom[ 1821]='h00000000;
    rd_cycle[ 1822] = 1'b0;  wr_cycle[ 1822] = 1'b1;  addr_rom[ 1822]='h00000474;  wr_data_rom[ 1822]='h00000543;
    rd_cycle[ 1823] = 1'b0;  wr_cycle[ 1823] = 1'b1;  addr_rom[ 1823]='h0000026c;  wr_data_rom[ 1823]='h000002e7;
    rd_cycle[ 1824] = 1'b0;  wr_cycle[ 1824] = 1'b1;  addr_rom[ 1824]='h000004e8;  wr_data_rom[ 1824]='h00000776;
    rd_cycle[ 1825] = 1'b0;  wr_cycle[ 1825] = 1'b1;  addr_rom[ 1825]='h00000444;  wr_data_rom[ 1825]='h0000057d;
    rd_cycle[ 1826] = 1'b0;  wr_cycle[ 1826] = 1'b1;  addr_rom[ 1826]='h000004a4;  wr_data_rom[ 1826]='h0000063d;
    rd_cycle[ 1827] = 1'b1;  wr_cycle[ 1827] = 1'b0;  addr_rom[ 1827]='h0000035c;  wr_data_rom[ 1827]='h00000000;
    rd_cycle[ 1828] = 1'b1;  wr_cycle[ 1828] = 1'b0;  addr_rom[ 1828]='h00000168;  wr_data_rom[ 1828]='h00000000;
    rd_cycle[ 1829] = 1'b0;  wr_cycle[ 1829] = 1'b1;  addr_rom[ 1829]='h0000004c;  wr_data_rom[ 1829]='h0000042c;
    rd_cycle[ 1830] = 1'b0;  wr_cycle[ 1830] = 1'b1;  addr_rom[ 1830]='h0000027c;  wr_data_rom[ 1830]='h000001e1;
    rd_cycle[ 1831] = 1'b0;  wr_cycle[ 1831] = 1'b1;  addr_rom[ 1831]='h0000004c;  wr_data_rom[ 1831]='h000003e1;
    rd_cycle[ 1832] = 1'b0;  wr_cycle[ 1832] = 1'b1;  addr_rom[ 1832]='h0000072c;  wr_data_rom[ 1832]='h0000027a;
    rd_cycle[ 1833] = 1'b1;  wr_cycle[ 1833] = 1'b0;  addr_rom[ 1833]='h00000034;  wr_data_rom[ 1833]='h00000000;
    rd_cycle[ 1834] = 1'b0;  wr_cycle[ 1834] = 1'b1;  addr_rom[ 1834]='h00000670;  wr_data_rom[ 1834]='h0000025f;
    rd_cycle[ 1835] = 1'b0;  wr_cycle[ 1835] = 1'b1;  addr_rom[ 1835]='h0000035c;  wr_data_rom[ 1835]='h000007e1;
    rd_cycle[ 1836] = 1'b0;  wr_cycle[ 1836] = 1'b1;  addr_rom[ 1836]='h000001d4;  wr_data_rom[ 1836]='h00000488;
    rd_cycle[ 1837] = 1'b1;  wr_cycle[ 1837] = 1'b0;  addr_rom[ 1837]='h0000052c;  wr_data_rom[ 1837]='h00000000;
    rd_cycle[ 1838] = 1'b1;  wr_cycle[ 1838] = 1'b0;  addr_rom[ 1838]='h00000388;  wr_data_rom[ 1838]='h00000000;
    rd_cycle[ 1839] = 1'b1;  wr_cycle[ 1839] = 1'b0;  addr_rom[ 1839]='h000006b8;  wr_data_rom[ 1839]='h00000000;
    rd_cycle[ 1840] = 1'b0;  wr_cycle[ 1840] = 1'b1;  addr_rom[ 1840]='h00000640;  wr_data_rom[ 1840]='h0000011f;
    rd_cycle[ 1841] = 1'b1;  wr_cycle[ 1841] = 1'b0;  addr_rom[ 1841]='h000001bc;  wr_data_rom[ 1841]='h00000000;
    rd_cycle[ 1842] = 1'b1;  wr_cycle[ 1842] = 1'b0;  addr_rom[ 1842]='h00000534;  wr_data_rom[ 1842]='h00000000;
    rd_cycle[ 1843] = 1'b0;  wr_cycle[ 1843] = 1'b1;  addr_rom[ 1843]='h0000065c;  wr_data_rom[ 1843]='h00000248;
    rd_cycle[ 1844] = 1'b0;  wr_cycle[ 1844] = 1'b1;  addr_rom[ 1844]='h00000048;  wr_data_rom[ 1844]='h00000578;
    rd_cycle[ 1845] = 1'b1;  wr_cycle[ 1845] = 1'b0;  addr_rom[ 1845]='h000004b0;  wr_data_rom[ 1845]='h00000000;
    rd_cycle[ 1846] = 1'b1;  wr_cycle[ 1846] = 1'b0;  addr_rom[ 1846]='h00000184;  wr_data_rom[ 1846]='h00000000;
    rd_cycle[ 1847] = 1'b1;  wr_cycle[ 1847] = 1'b0;  addr_rom[ 1847]='h0000072c;  wr_data_rom[ 1847]='h00000000;
    rd_cycle[ 1848] = 1'b1;  wr_cycle[ 1848] = 1'b0;  addr_rom[ 1848]='h00000004;  wr_data_rom[ 1848]='h00000000;
    rd_cycle[ 1849] = 1'b0;  wr_cycle[ 1849] = 1'b1;  addr_rom[ 1849]='h0000006c;  wr_data_rom[ 1849]='h000006c4;
    rd_cycle[ 1850] = 1'b1;  wr_cycle[ 1850] = 1'b0;  addr_rom[ 1850]='h000001f0;  wr_data_rom[ 1850]='h00000000;
    rd_cycle[ 1851] = 1'b0;  wr_cycle[ 1851] = 1'b1;  addr_rom[ 1851]='h00000420;  wr_data_rom[ 1851]='h00000595;
    rd_cycle[ 1852] = 1'b1;  wr_cycle[ 1852] = 1'b0;  addr_rom[ 1852]='h00000328;  wr_data_rom[ 1852]='h00000000;
    rd_cycle[ 1853] = 1'b1;  wr_cycle[ 1853] = 1'b0;  addr_rom[ 1853]='h00000630;  wr_data_rom[ 1853]='h00000000;
    rd_cycle[ 1854] = 1'b1;  wr_cycle[ 1854] = 1'b0;  addr_rom[ 1854]='h00000754;  wr_data_rom[ 1854]='h00000000;
    rd_cycle[ 1855] = 1'b0;  wr_cycle[ 1855] = 1'b1;  addr_rom[ 1855]='h0000031c;  wr_data_rom[ 1855]='h00000546;
    rd_cycle[ 1856] = 1'b1;  wr_cycle[ 1856] = 1'b0;  addr_rom[ 1856]='h00000430;  wr_data_rom[ 1856]='h00000000;
    rd_cycle[ 1857] = 1'b0;  wr_cycle[ 1857] = 1'b1;  addr_rom[ 1857]='h000003fc;  wr_data_rom[ 1857]='h000005b7;
    rd_cycle[ 1858] = 1'b1;  wr_cycle[ 1858] = 1'b0;  addr_rom[ 1858]='h0000077c;  wr_data_rom[ 1858]='h00000000;
    rd_cycle[ 1859] = 1'b0;  wr_cycle[ 1859] = 1'b1;  addr_rom[ 1859]='h00000324;  wr_data_rom[ 1859]='h000005e8;
    rd_cycle[ 1860] = 1'b1;  wr_cycle[ 1860] = 1'b0;  addr_rom[ 1860]='h000001b0;  wr_data_rom[ 1860]='h00000000;
    rd_cycle[ 1861] = 1'b0;  wr_cycle[ 1861] = 1'b1;  addr_rom[ 1861]='h000001c4;  wr_data_rom[ 1861]='h000003b4;
    rd_cycle[ 1862] = 1'b1;  wr_cycle[ 1862] = 1'b0;  addr_rom[ 1862]='h000005d0;  wr_data_rom[ 1862]='h00000000;
    rd_cycle[ 1863] = 1'b1;  wr_cycle[ 1863] = 1'b0;  addr_rom[ 1863]='h000001d4;  wr_data_rom[ 1863]='h00000000;
    rd_cycle[ 1864] = 1'b0;  wr_cycle[ 1864] = 1'b1;  addr_rom[ 1864]='h000006d8;  wr_data_rom[ 1864]='h000003e1;
    rd_cycle[ 1865] = 1'b0;  wr_cycle[ 1865] = 1'b1;  addr_rom[ 1865]='h00000114;  wr_data_rom[ 1865]='h00000316;
    rd_cycle[ 1866] = 1'b1;  wr_cycle[ 1866] = 1'b0;  addr_rom[ 1866]='h000005cc;  wr_data_rom[ 1866]='h00000000;
    rd_cycle[ 1867] = 1'b0;  wr_cycle[ 1867] = 1'b1;  addr_rom[ 1867]='h00000528;  wr_data_rom[ 1867]='h00000729;
    rd_cycle[ 1868] = 1'b0;  wr_cycle[ 1868] = 1'b1;  addr_rom[ 1868]='h00000054;  wr_data_rom[ 1868]='h00000377;
    rd_cycle[ 1869] = 1'b0;  wr_cycle[ 1869] = 1'b1;  addr_rom[ 1869]='h00000788;  wr_data_rom[ 1869]='h000000d1;
    rd_cycle[ 1870] = 1'b0;  wr_cycle[ 1870] = 1'b1;  addr_rom[ 1870]='h00000710;  wr_data_rom[ 1870]='h00000092;
    rd_cycle[ 1871] = 1'b1;  wr_cycle[ 1871] = 1'b0;  addr_rom[ 1871]='h0000017c;  wr_data_rom[ 1871]='h00000000;
    rd_cycle[ 1872] = 1'b0;  wr_cycle[ 1872] = 1'b1;  addr_rom[ 1872]='h00000194;  wr_data_rom[ 1872]='h0000015b;
    rd_cycle[ 1873] = 1'b1;  wr_cycle[ 1873] = 1'b0;  addr_rom[ 1873]='h000007f8;  wr_data_rom[ 1873]='h00000000;
    rd_cycle[ 1874] = 1'b1;  wr_cycle[ 1874] = 1'b0;  addr_rom[ 1874]='h0000024c;  wr_data_rom[ 1874]='h00000000;
    rd_cycle[ 1875] = 1'b1;  wr_cycle[ 1875] = 1'b0;  addr_rom[ 1875]='h00000080;  wr_data_rom[ 1875]='h00000000;
    rd_cycle[ 1876] = 1'b1;  wr_cycle[ 1876] = 1'b0;  addr_rom[ 1876]='h00000508;  wr_data_rom[ 1876]='h00000000;
    rd_cycle[ 1877] = 1'b0;  wr_cycle[ 1877] = 1'b1;  addr_rom[ 1877]='h000003a4;  wr_data_rom[ 1877]='h00000343;
    rd_cycle[ 1878] = 1'b0;  wr_cycle[ 1878] = 1'b1;  addr_rom[ 1878]='h0000048c;  wr_data_rom[ 1878]='h000006a9;
    rd_cycle[ 1879] = 1'b1;  wr_cycle[ 1879] = 1'b0;  addr_rom[ 1879]='h000000ec;  wr_data_rom[ 1879]='h00000000;
    rd_cycle[ 1880] = 1'b0;  wr_cycle[ 1880] = 1'b1;  addr_rom[ 1880]='h00000170;  wr_data_rom[ 1880]='h000004c0;
    rd_cycle[ 1881] = 1'b1;  wr_cycle[ 1881] = 1'b0;  addr_rom[ 1881]='h00000664;  wr_data_rom[ 1881]='h00000000;
    rd_cycle[ 1882] = 1'b1;  wr_cycle[ 1882] = 1'b0;  addr_rom[ 1882]='h000007ec;  wr_data_rom[ 1882]='h00000000;
    rd_cycle[ 1883] = 1'b1;  wr_cycle[ 1883] = 1'b0;  addr_rom[ 1883]='h00000778;  wr_data_rom[ 1883]='h00000000;
    rd_cycle[ 1884] = 1'b1;  wr_cycle[ 1884] = 1'b0;  addr_rom[ 1884]='h000001bc;  wr_data_rom[ 1884]='h00000000;
    rd_cycle[ 1885] = 1'b0;  wr_cycle[ 1885] = 1'b1;  addr_rom[ 1885]='h00000020;  wr_data_rom[ 1885]='h00000628;
    rd_cycle[ 1886] = 1'b0;  wr_cycle[ 1886] = 1'b1;  addr_rom[ 1886]='h00000094;  wr_data_rom[ 1886]='h00000547;
    rd_cycle[ 1887] = 1'b1;  wr_cycle[ 1887] = 1'b0;  addr_rom[ 1887]='h00000438;  wr_data_rom[ 1887]='h00000000;
    rd_cycle[ 1888] = 1'b1;  wr_cycle[ 1888] = 1'b0;  addr_rom[ 1888]='h000006b0;  wr_data_rom[ 1888]='h00000000;
    rd_cycle[ 1889] = 1'b1;  wr_cycle[ 1889] = 1'b0;  addr_rom[ 1889]='h00000544;  wr_data_rom[ 1889]='h00000000;
    rd_cycle[ 1890] = 1'b1;  wr_cycle[ 1890] = 1'b0;  addr_rom[ 1890]='h00000078;  wr_data_rom[ 1890]='h00000000;
    rd_cycle[ 1891] = 1'b0;  wr_cycle[ 1891] = 1'b1;  addr_rom[ 1891]='h0000032c;  wr_data_rom[ 1891]='h00000235;
    rd_cycle[ 1892] = 1'b0;  wr_cycle[ 1892] = 1'b1;  addr_rom[ 1892]='h00000300;  wr_data_rom[ 1892]='h0000033e;
    rd_cycle[ 1893] = 1'b0;  wr_cycle[ 1893] = 1'b1;  addr_rom[ 1893]='h00000550;  wr_data_rom[ 1893]='h000003cb;
    rd_cycle[ 1894] = 1'b0;  wr_cycle[ 1894] = 1'b1;  addr_rom[ 1894]='h000007ac;  wr_data_rom[ 1894]='h000001fc;
    rd_cycle[ 1895] = 1'b0;  wr_cycle[ 1895] = 1'b1;  addr_rom[ 1895]='h0000044c;  wr_data_rom[ 1895]='h0000076c;
    rd_cycle[ 1896] = 1'b1;  wr_cycle[ 1896] = 1'b0;  addr_rom[ 1896]='h000003d8;  wr_data_rom[ 1896]='h00000000;
    rd_cycle[ 1897] = 1'b1;  wr_cycle[ 1897] = 1'b0;  addr_rom[ 1897]='h00000354;  wr_data_rom[ 1897]='h00000000;
    rd_cycle[ 1898] = 1'b0;  wr_cycle[ 1898] = 1'b1;  addr_rom[ 1898]='h00000374;  wr_data_rom[ 1898]='h00000244;
    rd_cycle[ 1899] = 1'b0;  wr_cycle[ 1899] = 1'b1;  addr_rom[ 1899]='h00000130;  wr_data_rom[ 1899]='h00000002;
    rd_cycle[ 1900] = 1'b1;  wr_cycle[ 1900] = 1'b0;  addr_rom[ 1900]='h000007b4;  wr_data_rom[ 1900]='h00000000;
    rd_cycle[ 1901] = 1'b0;  wr_cycle[ 1901] = 1'b1;  addr_rom[ 1901]='h00000654;  wr_data_rom[ 1901]='h000004ec;
    rd_cycle[ 1902] = 1'b0;  wr_cycle[ 1902] = 1'b1;  addr_rom[ 1902]='h00000380;  wr_data_rom[ 1902]='h00000100;
    rd_cycle[ 1903] = 1'b1;  wr_cycle[ 1903] = 1'b0;  addr_rom[ 1903]='h000000d4;  wr_data_rom[ 1903]='h00000000;
    rd_cycle[ 1904] = 1'b1;  wr_cycle[ 1904] = 1'b0;  addr_rom[ 1904]='h00000188;  wr_data_rom[ 1904]='h00000000;
    rd_cycle[ 1905] = 1'b1;  wr_cycle[ 1905] = 1'b0;  addr_rom[ 1905]='h0000068c;  wr_data_rom[ 1905]='h00000000;
    rd_cycle[ 1906] = 1'b0;  wr_cycle[ 1906] = 1'b1;  addr_rom[ 1906]='h000005d0;  wr_data_rom[ 1906]='h00000705;
    rd_cycle[ 1907] = 1'b0;  wr_cycle[ 1907] = 1'b1;  addr_rom[ 1907]='h000005f4;  wr_data_rom[ 1907]='h000001b0;
    rd_cycle[ 1908] = 1'b0;  wr_cycle[ 1908] = 1'b1;  addr_rom[ 1908]='h00000108;  wr_data_rom[ 1908]='h00000406;
    rd_cycle[ 1909] = 1'b1;  wr_cycle[ 1909] = 1'b0;  addr_rom[ 1909]='h00000558;  wr_data_rom[ 1909]='h00000000;
    rd_cycle[ 1910] = 1'b1;  wr_cycle[ 1910] = 1'b0;  addr_rom[ 1910]='h000005d0;  wr_data_rom[ 1910]='h00000000;
    rd_cycle[ 1911] = 1'b1;  wr_cycle[ 1911] = 1'b0;  addr_rom[ 1911]='h000003c0;  wr_data_rom[ 1911]='h00000000;
    rd_cycle[ 1912] = 1'b0;  wr_cycle[ 1912] = 1'b1;  addr_rom[ 1912]='h00000264;  wr_data_rom[ 1912]='h000001c6;
    rd_cycle[ 1913] = 1'b1;  wr_cycle[ 1913] = 1'b0;  addr_rom[ 1913]='h000000a0;  wr_data_rom[ 1913]='h00000000;
    rd_cycle[ 1914] = 1'b0;  wr_cycle[ 1914] = 1'b1;  addr_rom[ 1914]='h000003d0;  wr_data_rom[ 1914]='h000004d6;
    rd_cycle[ 1915] = 1'b1;  wr_cycle[ 1915] = 1'b0;  addr_rom[ 1915]='h000004d4;  wr_data_rom[ 1915]='h00000000;
    rd_cycle[ 1916] = 1'b1;  wr_cycle[ 1916] = 1'b0;  addr_rom[ 1916]='h00000348;  wr_data_rom[ 1916]='h00000000;
    rd_cycle[ 1917] = 1'b0;  wr_cycle[ 1917] = 1'b1;  addr_rom[ 1917]='h00000218;  wr_data_rom[ 1917]='h000003ad;
    rd_cycle[ 1918] = 1'b0;  wr_cycle[ 1918] = 1'b1;  addr_rom[ 1918]='h000007bc;  wr_data_rom[ 1918]='h0000061e;
    rd_cycle[ 1919] = 1'b0;  wr_cycle[ 1919] = 1'b1;  addr_rom[ 1919]='h00000660;  wr_data_rom[ 1919]='h000001da;
    rd_cycle[ 1920] = 1'b0;  wr_cycle[ 1920] = 1'b1;  addr_rom[ 1920]='h0000003c;  wr_data_rom[ 1920]='h00000031;
    rd_cycle[ 1921] = 1'b1;  wr_cycle[ 1921] = 1'b0;  addr_rom[ 1921]='h00000490;  wr_data_rom[ 1921]='h00000000;
    rd_cycle[ 1922] = 1'b0;  wr_cycle[ 1922] = 1'b1;  addr_rom[ 1922]='h00000278;  wr_data_rom[ 1922]='h00000041;
    rd_cycle[ 1923] = 1'b1;  wr_cycle[ 1923] = 1'b0;  addr_rom[ 1923]='h000005d8;  wr_data_rom[ 1923]='h00000000;
    rd_cycle[ 1924] = 1'b1;  wr_cycle[ 1924] = 1'b0;  addr_rom[ 1924]='h0000054c;  wr_data_rom[ 1924]='h00000000;
    rd_cycle[ 1925] = 1'b0;  wr_cycle[ 1925] = 1'b1;  addr_rom[ 1925]='h000001fc;  wr_data_rom[ 1925]='h0000024f;
    rd_cycle[ 1926] = 1'b0;  wr_cycle[ 1926] = 1'b1;  addr_rom[ 1926]='h00000554;  wr_data_rom[ 1926]='h00000366;
    rd_cycle[ 1927] = 1'b1;  wr_cycle[ 1927] = 1'b0;  addr_rom[ 1927]='h00000330;  wr_data_rom[ 1927]='h00000000;
    rd_cycle[ 1928] = 1'b0;  wr_cycle[ 1928] = 1'b1;  addr_rom[ 1928]='h000007a0;  wr_data_rom[ 1928]='h00000175;
    rd_cycle[ 1929] = 1'b1;  wr_cycle[ 1929] = 1'b0;  addr_rom[ 1929]='h000006e0;  wr_data_rom[ 1929]='h00000000;
    rd_cycle[ 1930] = 1'b1;  wr_cycle[ 1930] = 1'b0;  addr_rom[ 1930]='h00000370;  wr_data_rom[ 1930]='h00000000;
    rd_cycle[ 1931] = 1'b1;  wr_cycle[ 1931] = 1'b0;  addr_rom[ 1931]='h00000680;  wr_data_rom[ 1931]='h00000000;
    rd_cycle[ 1932] = 1'b0;  wr_cycle[ 1932] = 1'b1;  addr_rom[ 1932]='h000004f0;  wr_data_rom[ 1932]='h000005f6;
    rd_cycle[ 1933] = 1'b1;  wr_cycle[ 1933] = 1'b0;  addr_rom[ 1933]='h0000059c;  wr_data_rom[ 1933]='h00000000;
    rd_cycle[ 1934] = 1'b0;  wr_cycle[ 1934] = 1'b1;  addr_rom[ 1934]='h00000458;  wr_data_rom[ 1934]='h00000489;
    rd_cycle[ 1935] = 1'b0;  wr_cycle[ 1935] = 1'b1;  addr_rom[ 1935]='h000007f8;  wr_data_rom[ 1935]='h000007e2;
    rd_cycle[ 1936] = 1'b1;  wr_cycle[ 1936] = 1'b0;  addr_rom[ 1936]='h000000e4;  wr_data_rom[ 1936]='h00000000;
    rd_cycle[ 1937] = 1'b0;  wr_cycle[ 1937] = 1'b1;  addr_rom[ 1937]='h000003bc;  wr_data_rom[ 1937]='h000002a5;
    rd_cycle[ 1938] = 1'b1;  wr_cycle[ 1938] = 1'b0;  addr_rom[ 1938]='h00000430;  wr_data_rom[ 1938]='h00000000;
    rd_cycle[ 1939] = 1'b1;  wr_cycle[ 1939] = 1'b0;  addr_rom[ 1939]='h00000184;  wr_data_rom[ 1939]='h00000000;
    rd_cycle[ 1940] = 1'b1;  wr_cycle[ 1940] = 1'b0;  addr_rom[ 1940]='h0000024c;  wr_data_rom[ 1940]='h00000000;
    rd_cycle[ 1941] = 1'b0;  wr_cycle[ 1941] = 1'b1;  addr_rom[ 1941]='h00000028;  wr_data_rom[ 1941]='h00000590;
    rd_cycle[ 1942] = 1'b0;  wr_cycle[ 1942] = 1'b1;  addr_rom[ 1942]='h0000057c;  wr_data_rom[ 1942]='h00000081;
    rd_cycle[ 1943] = 1'b0;  wr_cycle[ 1943] = 1'b1;  addr_rom[ 1943]='h0000037c;  wr_data_rom[ 1943]='h000005e4;
    rd_cycle[ 1944] = 1'b1;  wr_cycle[ 1944] = 1'b0;  addr_rom[ 1944]='h00000068;  wr_data_rom[ 1944]='h00000000;
    rd_cycle[ 1945] = 1'b0;  wr_cycle[ 1945] = 1'b1;  addr_rom[ 1945]='h0000059c;  wr_data_rom[ 1945]='h000002ea;
    rd_cycle[ 1946] = 1'b1;  wr_cycle[ 1946] = 1'b0;  addr_rom[ 1946]='h000003bc;  wr_data_rom[ 1946]='h00000000;
    rd_cycle[ 1947] = 1'b0;  wr_cycle[ 1947] = 1'b1;  addr_rom[ 1947]='h0000053c;  wr_data_rom[ 1947]='h000007e0;
    rd_cycle[ 1948] = 1'b1;  wr_cycle[ 1948] = 1'b0;  addr_rom[ 1948]='h000002a8;  wr_data_rom[ 1948]='h00000000;
    rd_cycle[ 1949] = 1'b1;  wr_cycle[ 1949] = 1'b0;  addr_rom[ 1949]='h00000384;  wr_data_rom[ 1949]='h00000000;
    rd_cycle[ 1950] = 1'b1;  wr_cycle[ 1950] = 1'b0;  addr_rom[ 1950]='h00000588;  wr_data_rom[ 1950]='h00000000;
    rd_cycle[ 1951] = 1'b0;  wr_cycle[ 1951] = 1'b1;  addr_rom[ 1951]='h000000f4;  wr_data_rom[ 1951]='h00000767;
    rd_cycle[ 1952] = 1'b0;  wr_cycle[ 1952] = 1'b1;  addr_rom[ 1952]='h00000430;  wr_data_rom[ 1952]='h00000068;
    rd_cycle[ 1953] = 1'b1;  wr_cycle[ 1953] = 1'b0;  addr_rom[ 1953]='h000002c8;  wr_data_rom[ 1953]='h00000000;
    rd_cycle[ 1954] = 1'b1;  wr_cycle[ 1954] = 1'b0;  addr_rom[ 1954]='h000005e8;  wr_data_rom[ 1954]='h00000000;
    rd_cycle[ 1955] = 1'b1;  wr_cycle[ 1955] = 1'b0;  addr_rom[ 1955]='h000002dc;  wr_data_rom[ 1955]='h00000000;
    rd_cycle[ 1956] = 1'b1;  wr_cycle[ 1956] = 1'b0;  addr_rom[ 1956]='h00000128;  wr_data_rom[ 1956]='h00000000;
    rd_cycle[ 1957] = 1'b0;  wr_cycle[ 1957] = 1'b1;  addr_rom[ 1957]='h00000458;  wr_data_rom[ 1957]='h00000153;
    rd_cycle[ 1958] = 1'b1;  wr_cycle[ 1958] = 1'b0;  addr_rom[ 1958]='h00000380;  wr_data_rom[ 1958]='h00000000;
    rd_cycle[ 1959] = 1'b0;  wr_cycle[ 1959] = 1'b1;  addr_rom[ 1959]='h00000474;  wr_data_rom[ 1959]='h00000024;
    rd_cycle[ 1960] = 1'b0;  wr_cycle[ 1960] = 1'b1;  addr_rom[ 1960]='h00000010;  wr_data_rom[ 1960]='h000006db;
    rd_cycle[ 1961] = 1'b0;  wr_cycle[ 1961] = 1'b1;  addr_rom[ 1961]='h00000070;  wr_data_rom[ 1961]='h0000036b;
    rd_cycle[ 1962] = 1'b1;  wr_cycle[ 1962] = 1'b0;  addr_rom[ 1962]='h000001b4;  wr_data_rom[ 1962]='h00000000;
    rd_cycle[ 1963] = 1'b0;  wr_cycle[ 1963] = 1'b1;  addr_rom[ 1963]='h000002d8;  wr_data_rom[ 1963]='h00000327;
    rd_cycle[ 1964] = 1'b0;  wr_cycle[ 1964] = 1'b1;  addr_rom[ 1964]='h000005c8;  wr_data_rom[ 1964]='h000007b9;
    rd_cycle[ 1965] = 1'b0;  wr_cycle[ 1965] = 1'b1;  addr_rom[ 1965]='h000003fc;  wr_data_rom[ 1965]='h00000223;
    rd_cycle[ 1966] = 1'b0;  wr_cycle[ 1966] = 1'b1;  addr_rom[ 1966]='h00000110;  wr_data_rom[ 1966]='h0000012f;
    rd_cycle[ 1967] = 1'b0;  wr_cycle[ 1967] = 1'b1;  addr_rom[ 1967]='h000006f4;  wr_data_rom[ 1967]='h00000605;
    rd_cycle[ 1968] = 1'b0;  wr_cycle[ 1968] = 1'b1;  addr_rom[ 1968]='h00000088;  wr_data_rom[ 1968]='h0000045a;
    rd_cycle[ 1969] = 1'b0;  wr_cycle[ 1969] = 1'b1;  addr_rom[ 1969]='h000003b8;  wr_data_rom[ 1969]='h00000587;
    rd_cycle[ 1970] = 1'b0;  wr_cycle[ 1970] = 1'b1;  addr_rom[ 1970]='h000000ac;  wr_data_rom[ 1970]='h00000536;
    rd_cycle[ 1971] = 1'b0;  wr_cycle[ 1971] = 1'b1;  addr_rom[ 1971]='h000005cc;  wr_data_rom[ 1971]='h000006a6;
    rd_cycle[ 1972] = 1'b0;  wr_cycle[ 1972] = 1'b1;  addr_rom[ 1972]='h00000260;  wr_data_rom[ 1972]='h000007d9;
    rd_cycle[ 1973] = 1'b1;  wr_cycle[ 1973] = 1'b0;  addr_rom[ 1973]='h0000013c;  wr_data_rom[ 1973]='h00000000;
    rd_cycle[ 1974] = 1'b0;  wr_cycle[ 1974] = 1'b1;  addr_rom[ 1974]='h000000ac;  wr_data_rom[ 1974]='h00000654;
    rd_cycle[ 1975] = 1'b1;  wr_cycle[ 1975] = 1'b0;  addr_rom[ 1975]='h00000638;  wr_data_rom[ 1975]='h00000000;
    rd_cycle[ 1976] = 1'b0;  wr_cycle[ 1976] = 1'b1;  addr_rom[ 1976]='h000006a4;  wr_data_rom[ 1976]='h0000040a;
    rd_cycle[ 1977] = 1'b0;  wr_cycle[ 1977] = 1'b1;  addr_rom[ 1977]='h000005e8;  wr_data_rom[ 1977]='h00000548;
    rd_cycle[ 1978] = 1'b1;  wr_cycle[ 1978] = 1'b0;  addr_rom[ 1978]='h00000208;  wr_data_rom[ 1978]='h00000000;
    rd_cycle[ 1979] = 1'b1;  wr_cycle[ 1979] = 1'b0;  addr_rom[ 1979]='h00000164;  wr_data_rom[ 1979]='h00000000;
    rd_cycle[ 1980] = 1'b0;  wr_cycle[ 1980] = 1'b1;  addr_rom[ 1980]='h00000310;  wr_data_rom[ 1980]='h00000589;
    rd_cycle[ 1981] = 1'b0;  wr_cycle[ 1981] = 1'b1;  addr_rom[ 1981]='h00000528;  wr_data_rom[ 1981]='h000000e4;
    rd_cycle[ 1982] = 1'b0;  wr_cycle[ 1982] = 1'b1;  addr_rom[ 1982]='h00000004;  wr_data_rom[ 1982]='h000006c4;
    rd_cycle[ 1983] = 1'b0;  wr_cycle[ 1983] = 1'b1;  addr_rom[ 1983]='h000003e8;  wr_data_rom[ 1983]='h00000224;
    rd_cycle[ 1984] = 1'b0;  wr_cycle[ 1984] = 1'b1;  addr_rom[ 1984]='h000005d8;  wr_data_rom[ 1984]='h000000a3;
    rd_cycle[ 1985] = 1'b1;  wr_cycle[ 1985] = 1'b0;  addr_rom[ 1985]='h00000438;  wr_data_rom[ 1985]='h00000000;
    rd_cycle[ 1986] = 1'b0;  wr_cycle[ 1986] = 1'b1;  addr_rom[ 1986]='h00000650;  wr_data_rom[ 1986]='h0000008c;
    rd_cycle[ 1987] = 1'b0;  wr_cycle[ 1987] = 1'b1;  addr_rom[ 1987]='h000004fc;  wr_data_rom[ 1987]='h000004a9;
    rd_cycle[ 1988] = 1'b1;  wr_cycle[ 1988] = 1'b0;  addr_rom[ 1988]='h00000558;  wr_data_rom[ 1988]='h00000000;
    rd_cycle[ 1989] = 1'b1;  wr_cycle[ 1989] = 1'b0;  addr_rom[ 1989]='h000007c4;  wr_data_rom[ 1989]='h00000000;
    rd_cycle[ 1990] = 1'b1;  wr_cycle[ 1990] = 1'b0;  addr_rom[ 1990]='h0000033c;  wr_data_rom[ 1990]='h00000000;
    rd_cycle[ 1991] = 1'b1;  wr_cycle[ 1991] = 1'b0;  addr_rom[ 1991]='h000002d8;  wr_data_rom[ 1991]='h00000000;
    rd_cycle[ 1992] = 1'b1;  wr_cycle[ 1992] = 1'b0;  addr_rom[ 1992]='h000001f8;  wr_data_rom[ 1992]='h00000000;
    rd_cycle[ 1993] = 1'b0;  wr_cycle[ 1993] = 1'b1;  addr_rom[ 1993]='h00000568;  wr_data_rom[ 1993]='h0000017b;
    rd_cycle[ 1994] = 1'b0;  wr_cycle[ 1994] = 1'b1;  addr_rom[ 1994]='h000001b4;  wr_data_rom[ 1994]='h0000022e;
    rd_cycle[ 1995] = 1'b0;  wr_cycle[ 1995] = 1'b1;  addr_rom[ 1995]='h00000708;  wr_data_rom[ 1995]='h0000050b;
    rd_cycle[ 1996] = 1'b1;  wr_cycle[ 1996] = 1'b0;  addr_rom[ 1996]='h000000c4;  wr_data_rom[ 1996]='h00000000;
    rd_cycle[ 1997] = 1'b1;  wr_cycle[ 1997] = 1'b0;  addr_rom[ 1997]='h00000394;  wr_data_rom[ 1997]='h00000000;
    rd_cycle[ 1998] = 1'b0;  wr_cycle[ 1998] = 1'b1;  addr_rom[ 1998]='h00000334;  wr_data_rom[ 1998]='h000002ba;
    rd_cycle[ 1999] = 1'b0;  wr_cycle[ 1999] = 1'b1;  addr_rom[ 1999]='h000005b8;  wr_data_rom[ 1999]='h00000339;
    rd_cycle[ 2000] = 1'b1;  wr_cycle[ 2000] = 1'b0;  addr_rom[ 2000]='h00000344;  wr_data_rom[ 2000]='h00000000;
    rd_cycle[ 2001] = 1'b0;  wr_cycle[ 2001] = 1'b1;  addr_rom[ 2001]='h0000067c;  wr_data_rom[ 2001]='h000006cd;
    rd_cycle[ 2002] = 1'b0;  wr_cycle[ 2002] = 1'b1;  addr_rom[ 2002]='h00000520;  wr_data_rom[ 2002]='h0000035b;
    rd_cycle[ 2003] = 1'b1;  wr_cycle[ 2003] = 1'b0;  addr_rom[ 2003]='h0000075c;  wr_data_rom[ 2003]='h00000000;
    rd_cycle[ 2004] = 1'b0;  wr_cycle[ 2004] = 1'b1;  addr_rom[ 2004]='h000004b0;  wr_data_rom[ 2004]='h000005a5;
    rd_cycle[ 2005] = 1'b0;  wr_cycle[ 2005] = 1'b1;  addr_rom[ 2005]='h0000056c;  wr_data_rom[ 2005]='h000007e9;
    rd_cycle[ 2006] = 1'b1;  wr_cycle[ 2006] = 1'b0;  addr_rom[ 2006]='h000007a4;  wr_data_rom[ 2006]='h00000000;
    rd_cycle[ 2007] = 1'b1;  wr_cycle[ 2007] = 1'b0;  addr_rom[ 2007]='h000007a4;  wr_data_rom[ 2007]='h00000000;
    rd_cycle[ 2008] = 1'b1;  wr_cycle[ 2008] = 1'b0;  addr_rom[ 2008]='h000003c8;  wr_data_rom[ 2008]='h00000000;
    rd_cycle[ 2009] = 1'b1;  wr_cycle[ 2009] = 1'b0;  addr_rom[ 2009]='h000006dc;  wr_data_rom[ 2009]='h00000000;
    rd_cycle[ 2010] = 1'b1;  wr_cycle[ 2010] = 1'b0;  addr_rom[ 2010]='h0000008c;  wr_data_rom[ 2010]='h00000000;
    rd_cycle[ 2011] = 1'b0;  wr_cycle[ 2011] = 1'b1;  addr_rom[ 2011]='h00000744;  wr_data_rom[ 2011]='h00000526;
    rd_cycle[ 2012] = 1'b1;  wr_cycle[ 2012] = 1'b0;  addr_rom[ 2012]='h0000000c;  wr_data_rom[ 2012]='h00000000;
    rd_cycle[ 2013] = 1'b0;  wr_cycle[ 2013] = 1'b1;  addr_rom[ 2013]='h000004d8;  wr_data_rom[ 2013]='h0000064e;
    rd_cycle[ 2014] = 1'b1;  wr_cycle[ 2014] = 1'b0;  addr_rom[ 2014]='h000007e4;  wr_data_rom[ 2014]='h00000000;
    rd_cycle[ 2015] = 1'b0;  wr_cycle[ 2015] = 1'b1;  addr_rom[ 2015]='h0000073c;  wr_data_rom[ 2015]='h000002eb;
    rd_cycle[ 2016] = 1'b1;  wr_cycle[ 2016] = 1'b0;  addr_rom[ 2016]='h00000214;  wr_data_rom[ 2016]='h00000000;
    rd_cycle[ 2017] = 1'b0;  wr_cycle[ 2017] = 1'b1;  addr_rom[ 2017]='h000002a8;  wr_data_rom[ 2017]='h0000059e;
    rd_cycle[ 2018] = 1'b0;  wr_cycle[ 2018] = 1'b1;  addr_rom[ 2018]='h00000380;  wr_data_rom[ 2018]='h00000597;
    rd_cycle[ 2019] = 1'b1;  wr_cycle[ 2019] = 1'b0;  addr_rom[ 2019]='h00000628;  wr_data_rom[ 2019]='h00000000;
    rd_cycle[ 2020] = 1'b0;  wr_cycle[ 2020] = 1'b1;  addr_rom[ 2020]='h00000608;  wr_data_rom[ 2020]='h0000056d;
    rd_cycle[ 2021] = 1'b0;  wr_cycle[ 2021] = 1'b1;  addr_rom[ 2021]='h000006d0;  wr_data_rom[ 2021]='h000000c3;
    rd_cycle[ 2022] = 1'b1;  wr_cycle[ 2022] = 1'b0;  addr_rom[ 2022]='h00000428;  wr_data_rom[ 2022]='h00000000;
    rd_cycle[ 2023] = 1'b0;  wr_cycle[ 2023] = 1'b1;  addr_rom[ 2023]='h000003a4;  wr_data_rom[ 2023]='h00000344;
    rd_cycle[ 2024] = 1'b1;  wr_cycle[ 2024] = 1'b0;  addr_rom[ 2024]='h00000038;  wr_data_rom[ 2024]='h00000000;
    rd_cycle[ 2025] = 1'b1;  wr_cycle[ 2025] = 1'b0;  addr_rom[ 2025]='h000001bc;  wr_data_rom[ 2025]='h00000000;
    rd_cycle[ 2026] = 1'b0;  wr_cycle[ 2026] = 1'b1;  addr_rom[ 2026]='h00000238;  wr_data_rom[ 2026]='h000003c9;
    rd_cycle[ 2027] = 1'b1;  wr_cycle[ 2027] = 1'b0;  addr_rom[ 2027]='h000001d4;  wr_data_rom[ 2027]='h00000000;
    rd_cycle[ 2028] = 1'b1;  wr_cycle[ 2028] = 1'b0;  addr_rom[ 2028]='h00000520;  wr_data_rom[ 2028]='h00000000;
    rd_cycle[ 2029] = 1'b0;  wr_cycle[ 2029] = 1'b1;  addr_rom[ 2029]='h0000001c;  wr_data_rom[ 2029]='h00000278;
    rd_cycle[ 2030] = 1'b1;  wr_cycle[ 2030] = 1'b0;  addr_rom[ 2030]='h0000012c;  wr_data_rom[ 2030]='h00000000;
    rd_cycle[ 2031] = 1'b1;  wr_cycle[ 2031] = 1'b0;  addr_rom[ 2031]='h00000244;  wr_data_rom[ 2031]='h00000000;
    rd_cycle[ 2032] = 1'b1;  wr_cycle[ 2032] = 1'b0;  addr_rom[ 2032]='h000006bc;  wr_data_rom[ 2032]='h00000000;
    rd_cycle[ 2033] = 1'b1;  wr_cycle[ 2033] = 1'b0;  addr_rom[ 2033]='h00000134;  wr_data_rom[ 2033]='h00000000;
    rd_cycle[ 2034] = 1'b0;  wr_cycle[ 2034] = 1'b1;  addr_rom[ 2034]='h0000067c;  wr_data_rom[ 2034]='h000005e0;
    rd_cycle[ 2035] = 1'b1;  wr_cycle[ 2035] = 1'b0;  addr_rom[ 2035]='h00000488;  wr_data_rom[ 2035]='h00000000;
    rd_cycle[ 2036] = 1'b0;  wr_cycle[ 2036] = 1'b1;  addr_rom[ 2036]='h00000510;  wr_data_rom[ 2036]='h000002a8;
    rd_cycle[ 2037] = 1'b1;  wr_cycle[ 2037] = 1'b0;  addr_rom[ 2037]='h000003c0;  wr_data_rom[ 2037]='h00000000;
    rd_cycle[ 2038] = 1'b0;  wr_cycle[ 2038] = 1'b1;  addr_rom[ 2038]='h000004a0;  wr_data_rom[ 2038]='h00000438;
    rd_cycle[ 2039] = 1'b0;  wr_cycle[ 2039] = 1'b1;  addr_rom[ 2039]='h00000704;  wr_data_rom[ 2039]='h00000527;
    rd_cycle[ 2040] = 1'b0;  wr_cycle[ 2040] = 1'b1;  addr_rom[ 2040]='h00000128;  wr_data_rom[ 2040]='h0000053f;
    rd_cycle[ 2041] = 1'b0;  wr_cycle[ 2041] = 1'b1;  addr_rom[ 2041]='h000001f4;  wr_data_rom[ 2041]='h0000074b;
    rd_cycle[ 2042] = 1'b1;  wr_cycle[ 2042] = 1'b0;  addr_rom[ 2042]='h00000684;  wr_data_rom[ 2042]='h00000000;
    rd_cycle[ 2043] = 1'b1;  wr_cycle[ 2043] = 1'b0;  addr_rom[ 2043]='h00000090;  wr_data_rom[ 2043]='h00000000;
    rd_cycle[ 2044] = 1'b1;  wr_cycle[ 2044] = 1'b0;  addr_rom[ 2044]='h00000728;  wr_data_rom[ 2044]='h00000000;
    rd_cycle[ 2045] = 1'b1;  wr_cycle[ 2045] = 1'b0;  addr_rom[ 2045]='h0000020c;  wr_data_rom[ 2045]='h00000000;
    rd_cycle[ 2046] = 1'b0;  wr_cycle[ 2046] = 1'b1;  addr_rom[ 2046]='h000002c4;  wr_data_rom[ 2046]='h00000555;
    rd_cycle[ 2047] = 1'b0;  wr_cycle[ 2047] = 1'b1;  addr_rom[ 2047]='h0000041c;  wr_data_rom[ 2047]='h000002ac;
    // 512 silence cycles
    rd_cycle[ 2048] = 1'b0;  wr_cycle[ 2048] = 1'b0;  addr_rom[ 2048]='h00000000;  wr_data_rom[ 2048]='h00000000;
    rd_cycle[ 2049] = 1'b0;  wr_cycle[ 2049] = 1'b0;  addr_rom[ 2049]='h00000000;  wr_data_rom[ 2049]='h00000000;
    rd_cycle[ 2050] = 1'b0;  wr_cycle[ 2050] = 1'b0;  addr_rom[ 2050]='h00000000;  wr_data_rom[ 2050]='h00000000;
    rd_cycle[ 2051] = 1'b0;  wr_cycle[ 2051] = 1'b0;  addr_rom[ 2051]='h00000000;  wr_data_rom[ 2051]='h00000000;
    rd_cycle[ 2052] = 1'b0;  wr_cycle[ 2052] = 1'b0;  addr_rom[ 2052]='h00000000;  wr_data_rom[ 2052]='h00000000;
    rd_cycle[ 2053] = 1'b0;  wr_cycle[ 2053] = 1'b0;  addr_rom[ 2053]='h00000000;  wr_data_rom[ 2053]='h00000000;
    rd_cycle[ 2054] = 1'b0;  wr_cycle[ 2054] = 1'b0;  addr_rom[ 2054]='h00000000;  wr_data_rom[ 2054]='h00000000;
    rd_cycle[ 2055] = 1'b0;  wr_cycle[ 2055] = 1'b0;  addr_rom[ 2055]='h00000000;  wr_data_rom[ 2055]='h00000000;
    rd_cycle[ 2056] = 1'b0;  wr_cycle[ 2056] = 1'b0;  addr_rom[ 2056]='h00000000;  wr_data_rom[ 2056]='h00000000;
    rd_cycle[ 2057] = 1'b0;  wr_cycle[ 2057] = 1'b0;  addr_rom[ 2057]='h00000000;  wr_data_rom[ 2057]='h00000000;
    rd_cycle[ 2058] = 1'b0;  wr_cycle[ 2058] = 1'b0;  addr_rom[ 2058]='h00000000;  wr_data_rom[ 2058]='h00000000;
    rd_cycle[ 2059] = 1'b0;  wr_cycle[ 2059] = 1'b0;  addr_rom[ 2059]='h00000000;  wr_data_rom[ 2059]='h00000000;
    rd_cycle[ 2060] = 1'b0;  wr_cycle[ 2060] = 1'b0;  addr_rom[ 2060]='h00000000;  wr_data_rom[ 2060]='h00000000;
    rd_cycle[ 2061] = 1'b0;  wr_cycle[ 2061] = 1'b0;  addr_rom[ 2061]='h00000000;  wr_data_rom[ 2061]='h00000000;
    rd_cycle[ 2062] = 1'b0;  wr_cycle[ 2062] = 1'b0;  addr_rom[ 2062]='h00000000;  wr_data_rom[ 2062]='h00000000;
    rd_cycle[ 2063] = 1'b0;  wr_cycle[ 2063] = 1'b0;  addr_rom[ 2063]='h00000000;  wr_data_rom[ 2063]='h00000000;
    rd_cycle[ 2064] = 1'b0;  wr_cycle[ 2064] = 1'b0;  addr_rom[ 2064]='h00000000;  wr_data_rom[ 2064]='h00000000;
    rd_cycle[ 2065] = 1'b0;  wr_cycle[ 2065] = 1'b0;  addr_rom[ 2065]='h00000000;  wr_data_rom[ 2065]='h00000000;
    rd_cycle[ 2066] = 1'b0;  wr_cycle[ 2066] = 1'b0;  addr_rom[ 2066]='h00000000;  wr_data_rom[ 2066]='h00000000;
    rd_cycle[ 2067] = 1'b0;  wr_cycle[ 2067] = 1'b0;  addr_rom[ 2067]='h00000000;  wr_data_rom[ 2067]='h00000000;
    rd_cycle[ 2068] = 1'b0;  wr_cycle[ 2068] = 1'b0;  addr_rom[ 2068]='h00000000;  wr_data_rom[ 2068]='h00000000;
    rd_cycle[ 2069] = 1'b0;  wr_cycle[ 2069] = 1'b0;  addr_rom[ 2069]='h00000000;  wr_data_rom[ 2069]='h00000000;
    rd_cycle[ 2070] = 1'b0;  wr_cycle[ 2070] = 1'b0;  addr_rom[ 2070]='h00000000;  wr_data_rom[ 2070]='h00000000;
    rd_cycle[ 2071] = 1'b0;  wr_cycle[ 2071] = 1'b0;  addr_rom[ 2071]='h00000000;  wr_data_rom[ 2071]='h00000000;
    rd_cycle[ 2072] = 1'b0;  wr_cycle[ 2072] = 1'b0;  addr_rom[ 2072]='h00000000;  wr_data_rom[ 2072]='h00000000;
    rd_cycle[ 2073] = 1'b0;  wr_cycle[ 2073] = 1'b0;  addr_rom[ 2073]='h00000000;  wr_data_rom[ 2073]='h00000000;
    rd_cycle[ 2074] = 1'b0;  wr_cycle[ 2074] = 1'b0;  addr_rom[ 2074]='h00000000;  wr_data_rom[ 2074]='h00000000;
    rd_cycle[ 2075] = 1'b0;  wr_cycle[ 2075] = 1'b0;  addr_rom[ 2075]='h00000000;  wr_data_rom[ 2075]='h00000000;
    rd_cycle[ 2076] = 1'b0;  wr_cycle[ 2076] = 1'b0;  addr_rom[ 2076]='h00000000;  wr_data_rom[ 2076]='h00000000;
    rd_cycle[ 2077] = 1'b0;  wr_cycle[ 2077] = 1'b0;  addr_rom[ 2077]='h00000000;  wr_data_rom[ 2077]='h00000000;
    rd_cycle[ 2078] = 1'b0;  wr_cycle[ 2078] = 1'b0;  addr_rom[ 2078]='h00000000;  wr_data_rom[ 2078]='h00000000;
    rd_cycle[ 2079] = 1'b0;  wr_cycle[ 2079] = 1'b0;  addr_rom[ 2079]='h00000000;  wr_data_rom[ 2079]='h00000000;
    rd_cycle[ 2080] = 1'b0;  wr_cycle[ 2080] = 1'b0;  addr_rom[ 2080]='h00000000;  wr_data_rom[ 2080]='h00000000;
    rd_cycle[ 2081] = 1'b0;  wr_cycle[ 2081] = 1'b0;  addr_rom[ 2081]='h00000000;  wr_data_rom[ 2081]='h00000000;
    rd_cycle[ 2082] = 1'b0;  wr_cycle[ 2082] = 1'b0;  addr_rom[ 2082]='h00000000;  wr_data_rom[ 2082]='h00000000;
    rd_cycle[ 2083] = 1'b0;  wr_cycle[ 2083] = 1'b0;  addr_rom[ 2083]='h00000000;  wr_data_rom[ 2083]='h00000000;
    rd_cycle[ 2084] = 1'b0;  wr_cycle[ 2084] = 1'b0;  addr_rom[ 2084]='h00000000;  wr_data_rom[ 2084]='h00000000;
    rd_cycle[ 2085] = 1'b0;  wr_cycle[ 2085] = 1'b0;  addr_rom[ 2085]='h00000000;  wr_data_rom[ 2085]='h00000000;
    rd_cycle[ 2086] = 1'b0;  wr_cycle[ 2086] = 1'b0;  addr_rom[ 2086]='h00000000;  wr_data_rom[ 2086]='h00000000;
    rd_cycle[ 2087] = 1'b0;  wr_cycle[ 2087] = 1'b0;  addr_rom[ 2087]='h00000000;  wr_data_rom[ 2087]='h00000000;
    rd_cycle[ 2088] = 1'b0;  wr_cycle[ 2088] = 1'b0;  addr_rom[ 2088]='h00000000;  wr_data_rom[ 2088]='h00000000;
    rd_cycle[ 2089] = 1'b0;  wr_cycle[ 2089] = 1'b0;  addr_rom[ 2089]='h00000000;  wr_data_rom[ 2089]='h00000000;
    rd_cycle[ 2090] = 1'b0;  wr_cycle[ 2090] = 1'b0;  addr_rom[ 2090]='h00000000;  wr_data_rom[ 2090]='h00000000;
    rd_cycle[ 2091] = 1'b0;  wr_cycle[ 2091] = 1'b0;  addr_rom[ 2091]='h00000000;  wr_data_rom[ 2091]='h00000000;
    rd_cycle[ 2092] = 1'b0;  wr_cycle[ 2092] = 1'b0;  addr_rom[ 2092]='h00000000;  wr_data_rom[ 2092]='h00000000;
    rd_cycle[ 2093] = 1'b0;  wr_cycle[ 2093] = 1'b0;  addr_rom[ 2093]='h00000000;  wr_data_rom[ 2093]='h00000000;
    rd_cycle[ 2094] = 1'b0;  wr_cycle[ 2094] = 1'b0;  addr_rom[ 2094]='h00000000;  wr_data_rom[ 2094]='h00000000;
    rd_cycle[ 2095] = 1'b0;  wr_cycle[ 2095] = 1'b0;  addr_rom[ 2095]='h00000000;  wr_data_rom[ 2095]='h00000000;
    rd_cycle[ 2096] = 1'b0;  wr_cycle[ 2096] = 1'b0;  addr_rom[ 2096]='h00000000;  wr_data_rom[ 2096]='h00000000;
    rd_cycle[ 2097] = 1'b0;  wr_cycle[ 2097] = 1'b0;  addr_rom[ 2097]='h00000000;  wr_data_rom[ 2097]='h00000000;
    rd_cycle[ 2098] = 1'b0;  wr_cycle[ 2098] = 1'b0;  addr_rom[ 2098]='h00000000;  wr_data_rom[ 2098]='h00000000;
    rd_cycle[ 2099] = 1'b0;  wr_cycle[ 2099] = 1'b0;  addr_rom[ 2099]='h00000000;  wr_data_rom[ 2099]='h00000000;
    rd_cycle[ 2100] = 1'b0;  wr_cycle[ 2100] = 1'b0;  addr_rom[ 2100]='h00000000;  wr_data_rom[ 2100]='h00000000;
    rd_cycle[ 2101] = 1'b0;  wr_cycle[ 2101] = 1'b0;  addr_rom[ 2101]='h00000000;  wr_data_rom[ 2101]='h00000000;
    rd_cycle[ 2102] = 1'b0;  wr_cycle[ 2102] = 1'b0;  addr_rom[ 2102]='h00000000;  wr_data_rom[ 2102]='h00000000;
    rd_cycle[ 2103] = 1'b0;  wr_cycle[ 2103] = 1'b0;  addr_rom[ 2103]='h00000000;  wr_data_rom[ 2103]='h00000000;
    rd_cycle[ 2104] = 1'b0;  wr_cycle[ 2104] = 1'b0;  addr_rom[ 2104]='h00000000;  wr_data_rom[ 2104]='h00000000;
    rd_cycle[ 2105] = 1'b0;  wr_cycle[ 2105] = 1'b0;  addr_rom[ 2105]='h00000000;  wr_data_rom[ 2105]='h00000000;
    rd_cycle[ 2106] = 1'b0;  wr_cycle[ 2106] = 1'b0;  addr_rom[ 2106]='h00000000;  wr_data_rom[ 2106]='h00000000;
    rd_cycle[ 2107] = 1'b0;  wr_cycle[ 2107] = 1'b0;  addr_rom[ 2107]='h00000000;  wr_data_rom[ 2107]='h00000000;
    rd_cycle[ 2108] = 1'b0;  wr_cycle[ 2108] = 1'b0;  addr_rom[ 2108]='h00000000;  wr_data_rom[ 2108]='h00000000;
    rd_cycle[ 2109] = 1'b0;  wr_cycle[ 2109] = 1'b0;  addr_rom[ 2109]='h00000000;  wr_data_rom[ 2109]='h00000000;
    rd_cycle[ 2110] = 1'b0;  wr_cycle[ 2110] = 1'b0;  addr_rom[ 2110]='h00000000;  wr_data_rom[ 2110]='h00000000;
    rd_cycle[ 2111] = 1'b0;  wr_cycle[ 2111] = 1'b0;  addr_rom[ 2111]='h00000000;  wr_data_rom[ 2111]='h00000000;
    rd_cycle[ 2112] = 1'b0;  wr_cycle[ 2112] = 1'b0;  addr_rom[ 2112]='h00000000;  wr_data_rom[ 2112]='h00000000;
    rd_cycle[ 2113] = 1'b0;  wr_cycle[ 2113] = 1'b0;  addr_rom[ 2113]='h00000000;  wr_data_rom[ 2113]='h00000000;
    rd_cycle[ 2114] = 1'b0;  wr_cycle[ 2114] = 1'b0;  addr_rom[ 2114]='h00000000;  wr_data_rom[ 2114]='h00000000;
    rd_cycle[ 2115] = 1'b0;  wr_cycle[ 2115] = 1'b0;  addr_rom[ 2115]='h00000000;  wr_data_rom[ 2115]='h00000000;
    rd_cycle[ 2116] = 1'b0;  wr_cycle[ 2116] = 1'b0;  addr_rom[ 2116]='h00000000;  wr_data_rom[ 2116]='h00000000;
    rd_cycle[ 2117] = 1'b0;  wr_cycle[ 2117] = 1'b0;  addr_rom[ 2117]='h00000000;  wr_data_rom[ 2117]='h00000000;
    rd_cycle[ 2118] = 1'b0;  wr_cycle[ 2118] = 1'b0;  addr_rom[ 2118]='h00000000;  wr_data_rom[ 2118]='h00000000;
    rd_cycle[ 2119] = 1'b0;  wr_cycle[ 2119] = 1'b0;  addr_rom[ 2119]='h00000000;  wr_data_rom[ 2119]='h00000000;
    rd_cycle[ 2120] = 1'b0;  wr_cycle[ 2120] = 1'b0;  addr_rom[ 2120]='h00000000;  wr_data_rom[ 2120]='h00000000;
    rd_cycle[ 2121] = 1'b0;  wr_cycle[ 2121] = 1'b0;  addr_rom[ 2121]='h00000000;  wr_data_rom[ 2121]='h00000000;
    rd_cycle[ 2122] = 1'b0;  wr_cycle[ 2122] = 1'b0;  addr_rom[ 2122]='h00000000;  wr_data_rom[ 2122]='h00000000;
    rd_cycle[ 2123] = 1'b0;  wr_cycle[ 2123] = 1'b0;  addr_rom[ 2123]='h00000000;  wr_data_rom[ 2123]='h00000000;
    rd_cycle[ 2124] = 1'b0;  wr_cycle[ 2124] = 1'b0;  addr_rom[ 2124]='h00000000;  wr_data_rom[ 2124]='h00000000;
    rd_cycle[ 2125] = 1'b0;  wr_cycle[ 2125] = 1'b0;  addr_rom[ 2125]='h00000000;  wr_data_rom[ 2125]='h00000000;
    rd_cycle[ 2126] = 1'b0;  wr_cycle[ 2126] = 1'b0;  addr_rom[ 2126]='h00000000;  wr_data_rom[ 2126]='h00000000;
    rd_cycle[ 2127] = 1'b0;  wr_cycle[ 2127] = 1'b0;  addr_rom[ 2127]='h00000000;  wr_data_rom[ 2127]='h00000000;
    rd_cycle[ 2128] = 1'b0;  wr_cycle[ 2128] = 1'b0;  addr_rom[ 2128]='h00000000;  wr_data_rom[ 2128]='h00000000;
    rd_cycle[ 2129] = 1'b0;  wr_cycle[ 2129] = 1'b0;  addr_rom[ 2129]='h00000000;  wr_data_rom[ 2129]='h00000000;
    rd_cycle[ 2130] = 1'b0;  wr_cycle[ 2130] = 1'b0;  addr_rom[ 2130]='h00000000;  wr_data_rom[ 2130]='h00000000;
    rd_cycle[ 2131] = 1'b0;  wr_cycle[ 2131] = 1'b0;  addr_rom[ 2131]='h00000000;  wr_data_rom[ 2131]='h00000000;
    rd_cycle[ 2132] = 1'b0;  wr_cycle[ 2132] = 1'b0;  addr_rom[ 2132]='h00000000;  wr_data_rom[ 2132]='h00000000;
    rd_cycle[ 2133] = 1'b0;  wr_cycle[ 2133] = 1'b0;  addr_rom[ 2133]='h00000000;  wr_data_rom[ 2133]='h00000000;
    rd_cycle[ 2134] = 1'b0;  wr_cycle[ 2134] = 1'b0;  addr_rom[ 2134]='h00000000;  wr_data_rom[ 2134]='h00000000;
    rd_cycle[ 2135] = 1'b0;  wr_cycle[ 2135] = 1'b0;  addr_rom[ 2135]='h00000000;  wr_data_rom[ 2135]='h00000000;
    rd_cycle[ 2136] = 1'b0;  wr_cycle[ 2136] = 1'b0;  addr_rom[ 2136]='h00000000;  wr_data_rom[ 2136]='h00000000;
    rd_cycle[ 2137] = 1'b0;  wr_cycle[ 2137] = 1'b0;  addr_rom[ 2137]='h00000000;  wr_data_rom[ 2137]='h00000000;
    rd_cycle[ 2138] = 1'b0;  wr_cycle[ 2138] = 1'b0;  addr_rom[ 2138]='h00000000;  wr_data_rom[ 2138]='h00000000;
    rd_cycle[ 2139] = 1'b0;  wr_cycle[ 2139] = 1'b0;  addr_rom[ 2139]='h00000000;  wr_data_rom[ 2139]='h00000000;
    rd_cycle[ 2140] = 1'b0;  wr_cycle[ 2140] = 1'b0;  addr_rom[ 2140]='h00000000;  wr_data_rom[ 2140]='h00000000;
    rd_cycle[ 2141] = 1'b0;  wr_cycle[ 2141] = 1'b0;  addr_rom[ 2141]='h00000000;  wr_data_rom[ 2141]='h00000000;
    rd_cycle[ 2142] = 1'b0;  wr_cycle[ 2142] = 1'b0;  addr_rom[ 2142]='h00000000;  wr_data_rom[ 2142]='h00000000;
    rd_cycle[ 2143] = 1'b0;  wr_cycle[ 2143] = 1'b0;  addr_rom[ 2143]='h00000000;  wr_data_rom[ 2143]='h00000000;
    rd_cycle[ 2144] = 1'b0;  wr_cycle[ 2144] = 1'b0;  addr_rom[ 2144]='h00000000;  wr_data_rom[ 2144]='h00000000;
    rd_cycle[ 2145] = 1'b0;  wr_cycle[ 2145] = 1'b0;  addr_rom[ 2145]='h00000000;  wr_data_rom[ 2145]='h00000000;
    rd_cycle[ 2146] = 1'b0;  wr_cycle[ 2146] = 1'b0;  addr_rom[ 2146]='h00000000;  wr_data_rom[ 2146]='h00000000;
    rd_cycle[ 2147] = 1'b0;  wr_cycle[ 2147] = 1'b0;  addr_rom[ 2147]='h00000000;  wr_data_rom[ 2147]='h00000000;
    rd_cycle[ 2148] = 1'b0;  wr_cycle[ 2148] = 1'b0;  addr_rom[ 2148]='h00000000;  wr_data_rom[ 2148]='h00000000;
    rd_cycle[ 2149] = 1'b0;  wr_cycle[ 2149] = 1'b0;  addr_rom[ 2149]='h00000000;  wr_data_rom[ 2149]='h00000000;
    rd_cycle[ 2150] = 1'b0;  wr_cycle[ 2150] = 1'b0;  addr_rom[ 2150]='h00000000;  wr_data_rom[ 2150]='h00000000;
    rd_cycle[ 2151] = 1'b0;  wr_cycle[ 2151] = 1'b0;  addr_rom[ 2151]='h00000000;  wr_data_rom[ 2151]='h00000000;
    rd_cycle[ 2152] = 1'b0;  wr_cycle[ 2152] = 1'b0;  addr_rom[ 2152]='h00000000;  wr_data_rom[ 2152]='h00000000;
    rd_cycle[ 2153] = 1'b0;  wr_cycle[ 2153] = 1'b0;  addr_rom[ 2153]='h00000000;  wr_data_rom[ 2153]='h00000000;
    rd_cycle[ 2154] = 1'b0;  wr_cycle[ 2154] = 1'b0;  addr_rom[ 2154]='h00000000;  wr_data_rom[ 2154]='h00000000;
    rd_cycle[ 2155] = 1'b0;  wr_cycle[ 2155] = 1'b0;  addr_rom[ 2155]='h00000000;  wr_data_rom[ 2155]='h00000000;
    rd_cycle[ 2156] = 1'b0;  wr_cycle[ 2156] = 1'b0;  addr_rom[ 2156]='h00000000;  wr_data_rom[ 2156]='h00000000;
    rd_cycle[ 2157] = 1'b0;  wr_cycle[ 2157] = 1'b0;  addr_rom[ 2157]='h00000000;  wr_data_rom[ 2157]='h00000000;
    rd_cycle[ 2158] = 1'b0;  wr_cycle[ 2158] = 1'b0;  addr_rom[ 2158]='h00000000;  wr_data_rom[ 2158]='h00000000;
    rd_cycle[ 2159] = 1'b0;  wr_cycle[ 2159] = 1'b0;  addr_rom[ 2159]='h00000000;  wr_data_rom[ 2159]='h00000000;
    rd_cycle[ 2160] = 1'b0;  wr_cycle[ 2160] = 1'b0;  addr_rom[ 2160]='h00000000;  wr_data_rom[ 2160]='h00000000;
    rd_cycle[ 2161] = 1'b0;  wr_cycle[ 2161] = 1'b0;  addr_rom[ 2161]='h00000000;  wr_data_rom[ 2161]='h00000000;
    rd_cycle[ 2162] = 1'b0;  wr_cycle[ 2162] = 1'b0;  addr_rom[ 2162]='h00000000;  wr_data_rom[ 2162]='h00000000;
    rd_cycle[ 2163] = 1'b0;  wr_cycle[ 2163] = 1'b0;  addr_rom[ 2163]='h00000000;  wr_data_rom[ 2163]='h00000000;
    rd_cycle[ 2164] = 1'b0;  wr_cycle[ 2164] = 1'b0;  addr_rom[ 2164]='h00000000;  wr_data_rom[ 2164]='h00000000;
    rd_cycle[ 2165] = 1'b0;  wr_cycle[ 2165] = 1'b0;  addr_rom[ 2165]='h00000000;  wr_data_rom[ 2165]='h00000000;
    rd_cycle[ 2166] = 1'b0;  wr_cycle[ 2166] = 1'b0;  addr_rom[ 2166]='h00000000;  wr_data_rom[ 2166]='h00000000;
    rd_cycle[ 2167] = 1'b0;  wr_cycle[ 2167] = 1'b0;  addr_rom[ 2167]='h00000000;  wr_data_rom[ 2167]='h00000000;
    rd_cycle[ 2168] = 1'b0;  wr_cycle[ 2168] = 1'b0;  addr_rom[ 2168]='h00000000;  wr_data_rom[ 2168]='h00000000;
    rd_cycle[ 2169] = 1'b0;  wr_cycle[ 2169] = 1'b0;  addr_rom[ 2169]='h00000000;  wr_data_rom[ 2169]='h00000000;
    rd_cycle[ 2170] = 1'b0;  wr_cycle[ 2170] = 1'b0;  addr_rom[ 2170]='h00000000;  wr_data_rom[ 2170]='h00000000;
    rd_cycle[ 2171] = 1'b0;  wr_cycle[ 2171] = 1'b0;  addr_rom[ 2171]='h00000000;  wr_data_rom[ 2171]='h00000000;
    rd_cycle[ 2172] = 1'b0;  wr_cycle[ 2172] = 1'b0;  addr_rom[ 2172]='h00000000;  wr_data_rom[ 2172]='h00000000;
    rd_cycle[ 2173] = 1'b0;  wr_cycle[ 2173] = 1'b0;  addr_rom[ 2173]='h00000000;  wr_data_rom[ 2173]='h00000000;
    rd_cycle[ 2174] = 1'b0;  wr_cycle[ 2174] = 1'b0;  addr_rom[ 2174]='h00000000;  wr_data_rom[ 2174]='h00000000;
    rd_cycle[ 2175] = 1'b0;  wr_cycle[ 2175] = 1'b0;  addr_rom[ 2175]='h00000000;  wr_data_rom[ 2175]='h00000000;
    rd_cycle[ 2176] = 1'b0;  wr_cycle[ 2176] = 1'b0;  addr_rom[ 2176]='h00000000;  wr_data_rom[ 2176]='h00000000;
    rd_cycle[ 2177] = 1'b0;  wr_cycle[ 2177] = 1'b0;  addr_rom[ 2177]='h00000000;  wr_data_rom[ 2177]='h00000000;
    rd_cycle[ 2178] = 1'b0;  wr_cycle[ 2178] = 1'b0;  addr_rom[ 2178]='h00000000;  wr_data_rom[ 2178]='h00000000;
    rd_cycle[ 2179] = 1'b0;  wr_cycle[ 2179] = 1'b0;  addr_rom[ 2179]='h00000000;  wr_data_rom[ 2179]='h00000000;
    rd_cycle[ 2180] = 1'b0;  wr_cycle[ 2180] = 1'b0;  addr_rom[ 2180]='h00000000;  wr_data_rom[ 2180]='h00000000;
    rd_cycle[ 2181] = 1'b0;  wr_cycle[ 2181] = 1'b0;  addr_rom[ 2181]='h00000000;  wr_data_rom[ 2181]='h00000000;
    rd_cycle[ 2182] = 1'b0;  wr_cycle[ 2182] = 1'b0;  addr_rom[ 2182]='h00000000;  wr_data_rom[ 2182]='h00000000;
    rd_cycle[ 2183] = 1'b0;  wr_cycle[ 2183] = 1'b0;  addr_rom[ 2183]='h00000000;  wr_data_rom[ 2183]='h00000000;
    rd_cycle[ 2184] = 1'b0;  wr_cycle[ 2184] = 1'b0;  addr_rom[ 2184]='h00000000;  wr_data_rom[ 2184]='h00000000;
    rd_cycle[ 2185] = 1'b0;  wr_cycle[ 2185] = 1'b0;  addr_rom[ 2185]='h00000000;  wr_data_rom[ 2185]='h00000000;
    rd_cycle[ 2186] = 1'b0;  wr_cycle[ 2186] = 1'b0;  addr_rom[ 2186]='h00000000;  wr_data_rom[ 2186]='h00000000;
    rd_cycle[ 2187] = 1'b0;  wr_cycle[ 2187] = 1'b0;  addr_rom[ 2187]='h00000000;  wr_data_rom[ 2187]='h00000000;
    rd_cycle[ 2188] = 1'b0;  wr_cycle[ 2188] = 1'b0;  addr_rom[ 2188]='h00000000;  wr_data_rom[ 2188]='h00000000;
    rd_cycle[ 2189] = 1'b0;  wr_cycle[ 2189] = 1'b0;  addr_rom[ 2189]='h00000000;  wr_data_rom[ 2189]='h00000000;
    rd_cycle[ 2190] = 1'b0;  wr_cycle[ 2190] = 1'b0;  addr_rom[ 2190]='h00000000;  wr_data_rom[ 2190]='h00000000;
    rd_cycle[ 2191] = 1'b0;  wr_cycle[ 2191] = 1'b0;  addr_rom[ 2191]='h00000000;  wr_data_rom[ 2191]='h00000000;
    rd_cycle[ 2192] = 1'b0;  wr_cycle[ 2192] = 1'b0;  addr_rom[ 2192]='h00000000;  wr_data_rom[ 2192]='h00000000;
    rd_cycle[ 2193] = 1'b0;  wr_cycle[ 2193] = 1'b0;  addr_rom[ 2193]='h00000000;  wr_data_rom[ 2193]='h00000000;
    rd_cycle[ 2194] = 1'b0;  wr_cycle[ 2194] = 1'b0;  addr_rom[ 2194]='h00000000;  wr_data_rom[ 2194]='h00000000;
    rd_cycle[ 2195] = 1'b0;  wr_cycle[ 2195] = 1'b0;  addr_rom[ 2195]='h00000000;  wr_data_rom[ 2195]='h00000000;
    rd_cycle[ 2196] = 1'b0;  wr_cycle[ 2196] = 1'b0;  addr_rom[ 2196]='h00000000;  wr_data_rom[ 2196]='h00000000;
    rd_cycle[ 2197] = 1'b0;  wr_cycle[ 2197] = 1'b0;  addr_rom[ 2197]='h00000000;  wr_data_rom[ 2197]='h00000000;
    rd_cycle[ 2198] = 1'b0;  wr_cycle[ 2198] = 1'b0;  addr_rom[ 2198]='h00000000;  wr_data_rom[ 2198]='h00000000;
    rd_cycle[ 2199] = 1'b0;  wr_cycle[ 2199] = 1'b0;  addr_rom[ 2199]='h00000000;  wr_data_rom[ 2199]='h00000000;
    rd_cycle[ 2200] = 1'b0;  wr_cycle[ 2200] = 1'b0;  addr_rom[ 2200]='h00000000;  wr_data_rom[ 2200]='h00000000;
    rd_cycle[ 2201] = 1'b0;  wr_cycle[ 2201] = 1'b0;  addr_rom[ 2201]='h00000000;  wr_data_rom[ 2201]='h00000000;
    rd_cycle[ 2202] = 1'b0;  wr_cycle[ 2202] = 1'b0;  addr_rom[ 2202]='h00000000;  wr_data_rom[ 2202]='h00000000;
    rd_cycle[ 2203] = 1'b0;  wr_cycle[ 2203] = 1'b0;  addr_rom[ 2203]='h00000000;  wr_data_rom[ 2203]='h00000000;
    rd_cycle[ 2204] = 1'b0;  wr_cycle[ 2204] = 1'b0;  addr_rom[ 2204]='h00000000;  wr_data_rom[ 2204]='h00000000;
    rd_cycle[ 2205] = 1'b0;  wr_cycle[ 2205] = 1'b0;  addr_rom[ 2205]='h00000000;  wr_data_rom[ 2205]='h00000000;
    rd_cycle[ 2206] = 1'b0;  wr_cycle[ 2206] = 1'b0;  addr_rom[ 2206]='h00000000;  wr_data_rom[ 2206]='h00000000;
    rd_cycle[ 2207] = 1'b0;  wr_cycle[ 2207] = 1'b0;  addr_rom[ 2207]='h00000000;  wr_data_rom[ 2207]='h00000000;
    rd_cycle[ 2208] = 1'b0;  wr_cycle[ 2208] = 1'b0;  addr_rom[ 2208]='h00000000;  wr_data_rom[ 2208]='h00000000;
    rd_cycle[ 2209] = 1'b0;  wr_cycle[ 2209] = 1'b0;  addr_rom[ 2209]='h00000000;  wr_data_rom[ 2209]='h00000000;
    rd_cycle[ 2210] = 1'b0;  wr_cycle[ 2210] = 1'b0;  addr_rom[ 2210]='h00000000;  wr_data_rom[ 2210]='h00000000;
    rd_cycle[ 2211] = 1'b0;  wr_cycle[ 2211] = 1'b0;  addr_rom[ 2211]='h00000000;  wr_data_rom[ 2211]='h00000000;
    rd_cycle[ 2212] = 1'b0;  wr_cycle[ 2212] = 1'b0;  addr_rom[ 2212]='h00000000;  wr_data_rom[ 2212]='h00000000;
    rd_cycle[ 2213] = 1'b0;  wr_cycle[ 2213] = 1'b0;  addr_rom[ 2213]='h00000000;  wr_data_rom[ 2213]='h00000000;
    rd_cycle[ 2214] = 1'b0;  wr_cycle[ 2214] = 1'b0;  addr_rom[ 2214]='h00000000;  wr_data_rom[ 2214]='h00000000;
    rd_cycle[ 2215] = 1'b0;  wr_cycle[ 2215] = 1'b0;  addr_rom[ 2215]='h00000000;  wr_data_rom[ 2215]='h00000000;
    rd_cycle[ 2216] = 1'b0;  wr_cycle[ 2216] = 1'b0;  addr_rom[ 2216]='h00000000;  wr_data_rom[ 2216]='h00000000;
    rd_cycle[ 2217] = 1'b0;  wr_cycle[ 2217] = 1'b0;  addr_rom[ 2217]='h00000000;  wr_data_rom[ 2217]='h00000000;
    rd_cycle[ 2218] = 1'b0;  wr_cycle[ 2218] = 1'b0;  addr_rom[ 2218]='h00000000;  wr_data_rom[ 2218]='h00000000;
    rd_cycle[ 2219] = 1'b0;  wr_cycle[ 2219] = 1'b0;  addr_rom[ 2219]='h00000000;  wr_data_rom[ 2219]='h00000000;
    rd_cycle[ 2220] = 1'b0;  wr_cycle[ 2220] = 1'b0;  addr_rom[ 2220]='h00000000;  wr_data_rom[ 2220]='h00000000;
    rd_cycle[ 2221] = 1'b0;  wr_cycle[ 2221] = 1'b0;  addr_rom[ 2221]='h00000000;  wr_data_rom[ 2221]='h00000000;
    rd_cycle[ 2222] = 1'b0;  wr_cycle[ 2222] = 1'b0;  addr_rom[ 2222]='h00000000;  wr_data_rom[ 2222]='h00000000;
    rd_cycle[ 2223] = 1'b0;  wr_cycle[ 2223] = 1'b0;  addr_rom[ 2223]='h00000000;  wr_data_rom[ 2223]='h00000000;
    rd_cycle[ 2224] = 1'b0;  wr_cycle[ 2224] = 1'b0;  addr_rom[ 2224]='h00000000;  wr_data_rom[ 2224]='h00000000;
    rd_cycle[ 2225] = 1'b0;  wr_cycle[ 2225] = 1'b0;  addr_rom[ 2225]='h00000000;  wr_data_rom[ 2225]='h00000000;
    rd_cycle[ 2226] = 1'b0;  wr_cycle[ 2226] = 1'b0;  addr_rom[ 2226]='h00000000;  wr_data_rom[ 2226]='h00000000;
    rd_cycle[ 2227] = 1'b0;  wr_cycle[ 2227] = 1'b0;  addr_rom[ 2227]='h00000000;  wr_data_rom[ 2227]='h00000000;
    rd_cycle[ 2228] = 1'b0;  wr_cycle[ 2228] = 1'b0;  addr_rom[ 2228]='h00000000;  wr_data_rom[ 2228]='h00000000;
    rd_cycle[ 2229] = 1'b0;  wr_cycle[ 2229] = 1'b0;  addr_rom[ 2229]='h00000000;  wr_data_rom[ 2229]='h00000000;
    rd_cycle[ 2230] = 1'b0;  wr_cycle[ 2230] = 1'b0;  addr_rom[ 2230]='h00000000;  wr_data_rom[ 2230]='h00000000;
    rd_cycle[ 2231] = 1'b0;  wr_cycle[ 2231] = 1'b0;  addr_rom[ 2231]='h00000000;  wr_data_rom[ 2231]='h00000000;
    rd_cycle[ 2232] = 1'b0;  wr_cycle[ 2232] = 1'b0;  addr_rom[ 2232]='h00000000;  wr_data_rom[ 2232]='h00000000;
    rd_cycle[ 2233] = 1'b0;  wr_cycle[ 2233] = 1'b0;  addr_rom[ 2233]='h00000000;  wr_data_rom[ 2233]='h00000000;
    rd_cycle[ 2234] = 1'b0;  wr_cycle[ 2234] = 1'b0;  addr_rom[ 2234]='h00000000;  wr_data_rom[ 2234]='h00000000;
    rd_cycle[ 2235] = 1'b0;  wr_cycle[ 2235] = 1'b0;  addr_rom[ 2235]='h00000000;  wr_data_rom[ 2235]='h00000000;
    rd_cycle[ 2236] = 1'b0;  wr_cycle[ 2236] = 1'b0;  addr_rom[ 2236]='h00000000;  wr_data_rom[ 2236]='h00000000;
    rd_cycle[ 2237] = 1'b0;  wr_cycle[ 2237] = 1'b0;  addr_rom[ 2237]='h00000000;  wr_data_rom[ 2237]='h00000000;
    rd_cycle[ 2238] = 1'b0;  wr_cycle[ 2238] = 1'b0;  addr_rom[ 2238]='h00000000;  wr_data_rom[ 2238]='h00000000;
    rd_cycle[ 2239] = 1'b0;  wr_cycle[ 2239] = 1'b0;  addr_rom[ 2239]='h00000000;  wr_data_rom[ 2239]='h00000000;
    rd_cycle[ 2240] = 1'b0;  wr_cycle[ 2240] = 1'b0;  addr_rom[ 2240]='h00000000;  wr_data_rom[ 2240]='h00000000;
    rd_cycle[ 2241] = 1'b0;  wr_cycle[ 2241] = 1'b0;  addr_rom[ 2241]='h00000000;  wr_data_rom[ 2241]='h00000000;
    rd_cycle[ 2242] = 1'b0;  wr_cycle[ 2242] = 1'b0;  addr_rom[ 2242]='h00000000;  wr_data_rom[ 2242]='h00000000;
    rd_cycle[ 2243] = 1'b0;  wr_cycle[ 2243] = 1'b0;  addr_rom[ 2243]='h00000000;  wr_data_rom[ 2243]='h00000000;
    rd_cycle[ 2244] = 1'b0;  wr_cycle[ 2244] = 1'b0;  addr_rom[ 2244]='h00000000;  wr_data_rom[ 2244]='h00000000;
    rd_cycle[ 2245] = 1'b0;  wr_cycle[ 2245] = 1'b0;  addr_rom[ 2245]='h00000000;  wr_data_rom[ 2245]='h00000000;
    rd_cycle[ 2246] = 1'b0;  wr_cycle[ 2246] = 1'b0;  addr_rom[ 2246]='h00000000;  wr_data_rom[ 2246]='h00000000;
    rd_cycle[ 2247] = 1'b0;  wr_cycle[ 2247] = 1'b0;  addr_rom[ 2247]='h00000000;  wr_data_rom[ 2247]='h00000000;
    rd_cycle[ 2248] = 1'b0;  wr_cycle[ 2248] = 1'b0;  addr_rom[ 2248]='h00000000;  wr_data_rom[ 2248]='h00000000;
    rd_cycle[ 2249] = 1'b0;  wr_cycle[ 2249] = 1'b0;  addr_rom[ 2249]='h00000000;  wr_data_rom[ 2249]='h00000000;
    rd_cycle[ 2250] = 1'b0;  wr_cycle[ 2250] = 1'b0;  addr_rom[ 2250]='h00000000;  wr_data_rom[ 2250]='h00000000;
    rd_cycle[ 2251] = 1'b0;  wr_cycle[ 2251] = 1'b0;  addr_rom[ 2251]='h00000000;  wr_data_rom[ 2251]='h00000000;
    rd_cycle[ 2252] = 1'b0;  wr_cycle[ 2252] = 1'b0;  addr_rom[ 2252]='h00000000;  wr_data_rom[ 2252]='h00000000;
    rd_cycle[ 2253] = 1'b0;  wr_cycle[ 2253] = 1'b0;  addr_rom[ 2253]='h00000000;  wr_data_rom[ 2253]='h00000000;
    rd_cycle[ 2254] = 1'b0;  wr_cycle[ 2254] = 1'b0;  addr_rom[ 2254]='h00000000;  wr_data_rom[ 2254]='h00000000;
    rd_cycle[ 2255] = 1'b0;  wr_cycle[ 2255] = 1'b0;  addr_rom[ 2255]='h00000000;  wr_data_rom[ 2255]='h00000000;
    rd_cycle[ 2256] = 1'b0;  wr_cycle[ 2256] = 1'b0;  addr_rom[ 2256]='h00000000;  wr_data_rom[ 2256]='h00000000;
    rd_cycle[ 2257] = 1'b0;  wr_cycle[ 2257] = 1'b0;  addr_rom[ 2257]='h00000000;  wr_data_rom[ 2257]='h00000000;
    rd_cycle[ 2258] = 1'b0;  wr_cycle[ 2258] = 1'b0;  addr_rom[ 2258]='h00000000;  wr_data_rom[ 2258]='h00000000;
    rd_cycle[ 2259] = 1'b0;  wr_cycle[ 2259] = 1'b0;  addr_rom[ 2259]='h00000000;  wr_data_rom[ 2259]='h00000000;
    rd_cycle[ 2260] = 1'b0;  wr_cycle[ 2260] = 1'b0;  addr_rom[ 2260]='h00000000;  wr_data_rom[ 2260]='h00000000;
    rd_cycle[ 2261] = 1'b0;  wr_cycle[ 2261] = 1'b0;  addr_rom[ 2261]='h00000000;  wr_data_rom[ 2261]='h00000000;
    rd_cycle[ 2262] = 1'b0;  wr_cycle[ 2262] = 1'b0;  addr_rom[ 2262]='h00000000;  wr_data_rom[ 2262]='h00000000;
    rd_cycle[ 2263] = 1'b0;  wr_cycle[ 2263] = 1'b0;  addr_rom[ 2263]='h00000000;  wr_data_rom[ 2263]='h00000000;
    rd_cycle[ 2264] = 1'b0;  wr_cycle[ 2264] = 1'b0;  addr_rom[ 2264]='h00000000;  wr_data_rom[ 2264]='h00000000;
    rd_cycle[ 2265] = 1'b0;  wr_cycle[ 2265] = 1'b0;  addr_rom[ 2265]='h00000000;  wr_data_rom[ 2265]='h00000000;
    rd_cycle[ 2266] = 1'b0;  wr_cycle[ 2266] = 1'b0;  addr_rom[ 2266]='h00000000;  wr_data_rom[ 2266]='h00000000;
    rd_cycle[ 2267] = 1'b0;  wr_cycle[ 2267] = 1'b0;  addr_rom[ 2267]='h00000000;  wr_data_rom[ 2267]='h00000000;
    rd_cycle[ 2268] = 1'b0;  wr_cycle[ 2268] = 1'b0;  addr_rom[ 2268]='h00000000;  wr_data_rom[ 2268]='h00000000;
    rd_cycle[ 2269] = 1'b0;  wr_cycle[ 2269] = 1'b0;  addr_rom[ 2269]='h00000000;  wr_data_rom[ 2269]='h00000000;
    rd_cycle[ 2270] = 1'b0;  wr_cycle[ 2270] = 1'b0;  addr_rom[ 2270]='h00000000;  wr_data_rom[ 2270]='h00000000;
    rd_cycle[ 2271] = 1'b0;  wr_cycle[ 2271] = 1'b0;  addr_rom[ 2271]='h00000000;  wr_data_rom[ 2271]='h00000000;
    rd_cycle[ 2272] = 1'b0;  wr_cycle[ 2272] = 1'b0;  addr_rom[ 2272]='h00000000;  wr_data_rom[ 2272]='h00000000;
    rd_cycle[ 2273] = 1'b0;  wr_cycle[ 2273] = 1'b0;  addr_rom[ 2273]='h00000000;  wr_data_rom[ 2273]='h00000000;
    rd_cycle[ 2274] = 1'b0;  wr_cycle[ 2274] = 1'b0;  addr_rom[ 2274]='h00000000;  wr_data_rom[ 2274]='h00000000;
    rd_cycle[ 2275] = 1'b0;  wr_cycle[ 2275] = 1'b0;  addr_rom[ 2275]='h00000000;  wr_data_rom[ 2275]='h00000000;
    rd_cycle[ 2276] = 1'b0;  wr_cycle[ 2276] = 1'b0;  addr_rom[ 2276]='h00000000;  wr_data_rom[ 2276]='h00000000;
    rd_cycle[ 2277] = 1'b0;  wr_cycle[ 2277] = 1'b0;  addr_rom[ 2277]='h00000000;  wr_data_rom[ 2277]='h00000000;
    rd_cycle[ 2278] = 1'b0;  wr_cycle[ 2278] = 1'b0;  addr_rom[ 2278]='h00000000;  wr_data_rom[ 2278]='h00000000;
    rd_cycle[ 2279] = 1'b0;  wr_cycle[ 2279] = 1'b0;  addr_rom[ 2279]='h00000000;  wr_data_rom[ 2279]='h00000000;
    rd_cycle[ 2280] = 1'b0;  wr_cycle[ 2280] = 1'b0;  addr_rom[ 2280]='h00000000;  wr_data_rom[ 2280]='h00000000;
    rd_cycle[ 2281] = 1'b0;  wr_cycle[ 2281] = 1'b0;  addr_rom[ 2281]='h00000000;  wr_data_rom[ 2281]='h00000000;
    rd_cycle[ 2282] = 1'b0;  wr_cycle[ 2282] = 1'b0;  addr_rom[ 2282]='h00000000;  wr_data_rom[ 2282]='h00000000;
    rd_cycle[ 2283] = 1'b0;  wr_cycle[ 2283] = 1'b0;  addr_rom[ 2283]='h00000000;  wr_data_rom[ 2283]='h00000000;
    rd_cycle[ 2284] = 1'b0;  wr_cycle[ 2284] = 1'b0;  addr_rom[ 2284]='h00000000;  wr_data_rom[ 2284]='h00000000;
    rd_cycle[ 2285] = 1'b0;  wr_cycle[ 2285] = 1'b0;  addr_rom[ 2285]='h00000000;  wr_data_rom[ 2285]='h00000000;
    rd_cycle[ 2286] = 1'b0;  wr_cycle[ 2286] = 1'b0;  addr_rom[ 2286]='h00000000;  wr_data_rom[ 2286]='h00000000;
    rd_cycle[ 2287] = 1'b0;  wr_cycle[ 2287] = 1'b0;  addr_rom[ 2287]='h00000000;  wr_data_rom[ 2287]='h00000000;
    rd_cycle[ 2288] = 1'b0;  wr_cycle[ 2288] = 1'b0;  addr_rom[ 2288]='h00000000;  wr_data_rom[ 2288]='h00000000;
    rd_cycle[ 2289] = 1'b0;  wr_cycle[ 2289] = 1'b0;  addr_rom[ 2289]='h00000000;  wr_data_rom[ 2289]='h00000000;
    rd_cycle[ 2290] = 1'b0;  wr_cycle[ 2290] = 1'b0;  addr_rom[ 2290]='h00000000;  wr_data_rom[ 2290]='h00000000;
    rd_cycle[ 2291] = 1'b0;  wr_cycle[ 2291] = 1'b0;  addr_rom[ 2291]='h00000000;  wr_data_rom[ 2291]='h00000000;
    rd_cycle[ 2292] = 1'b0;  wr_cycle[ 2292] = 1'b0;  addr_rom[ 2292]='h00000000;  wr_data_rom[ 2292]='h00000000;
    rd_cycle[ 2293] = 1'b0;  wr_cycle[ 2293] = 1'b0;  addr_rom[ 2293]='h00000000;  wr_data_rom[ 2293]='h00000000;
    rd_cycle[ 2294] = 1'b0;  wr_cycle[ 2294] = 1'b0;  addr_rom[ 2294]='h00000000;  wr_data_rom[ 2294]='h00000000;
    rd_cycle[ 2295] = 1'b0;  wr_cycle[ 2295] = 1'b0;  addr_rom[ 2295]='h00000000;  wr_data_rom[ 2295]='h00000000;
    rd_cycle[ 2296] = 1'b0;  wr_cycle[ 2296] = 1'b0;  addr_rom[ 2296]='h00000000;  wr_data_rom[ 2296]='h00000000;
    rd_cycle[ 2297] = 1'b0;  wr_cycle[ 2297] = 1'b0;  addr_rom[ 2297]='h00000000;  wr_data_rom[ 2297]='h00000000;
    rd_cycle[ 2298] = 1'b0;  wr_cycle[ 2298] = 1'b0;  addr_rom[ 2298]='h00000000;  wr_data_rom[ 2298]='h00000000;
    rd_cycle[ 2299] = 1'b0;  wr_cycle[ 2299] = 1'b0;  addr_rom[ 2299]='h00000000;  wr_data_rom[ 2299]='h00000000;
    rd_cycle[ 2300] = 1'b0;  wr_cycle[ 2300] = 1'b0;  addr_rom[ 2300]='h00000000;  wr_data_rom[ 2300]='h00000000;
    rd_cycle[ 2301] = 1'b0;  wr_cycle[ 2301] = 1'b0;  addr_rom[ 2301]='h00000000;  wr_data_rom[ 2301]='h00000000;
    rd_cycle[ 2302] = 1'b0;  wr_cycle[ 2302] = 1'b0;  addr_rom[ 2302]='h00000000;  wr_data_rom[ 2302]='h00000000;
    rd_cycle[ 2303] = 1'b0;  wr_cycle[ 2303] = 1'b0;  addr_rom[ 2303]='h00000000;  wr_data_rom[ 2303]='h00000000;
    rd_cycle[ 2304] = 1'b0;  wr_cycle[ 2304] = 1'b0;  addr_rom[ 2304]='h00000000;  wr_data_rom[ 2304]='h00000000;
    rd_cycle[ 2305] = 1'b0;  wr_cycle[ 2305] = 1'b0;  addr_rom[ 2305]='h00000000;  wr_data_rom[ 2305]='h00000000;
    rd_cycle[ 2306] = 1'b0;  wr_cycle[ 2306] = 1'b0;  addr_rom[ 2306]='h00000000;  wr_data_rom[ 2306]='h00000000;
    rd_cycle[ 2307] = 1'b0;  wr_cycle[ 2307] = 1'b0;  addr_rom[ 2307]='h00000000;  wr_data_rom[ 2307]='h00000000;
    rd_cycle[ 2308] = 1'b0;  wr_cycle[ 2308] = 1'b0;  addr_rom[ 2308]='h00000000;  wr_data_rom[ 2308]='h00000000;
    rd_cycle[ 2309] = 1'b0;  wr_cycle[ 2309] = 1'b0;  addr_rom[ 2309]='h00000000;  wr_data_rom[ 2309]='h00000000;
    rd_cycle[ 2310] = 1'b0;  wr_cycle[ 2310] = 1'b0;  addr_rom[ 2310]='h00000000;  wr_data_rom[ 2310]='h00000000;
    rd_cycle[ 2311] = 1'b0;  wr_cycle[ 2311] = 1'b0;  addr_rom[ 2311]='h00000000;  wr_data_rom[ 2311]='h00000000;
    rd_cycle[ 2312] = 1'b0;  wr_cycle[ 2312] = 1'b0;  addr_rom[ 2312]='h00000000;  wr_data_rom[ 2312]='h00000000;
    rd_cycle[ 2313] = 1'b0;  wr_cycle[ 2313] = 1'b0;  addr_rom[ 2313]='h00000000;  wr_data_rom[ 2313]='h00000000;
    rd_cycle[ 2314] = 1'b0;  wr_cycle[ 2314] = 1'b0;  addr_rom[ 2314]='h00000000;  wr_data_rom[ 2314]='h00000000;
    rd_cycle[ 2315] = 1'b0;  wr_cycle[ 2315] = 1'b0;  addr_rom[ 2315]='h00000000;  wr_data_rom[ 2315]='h00000000;
    rd_cycle[ 2316] = 1'b0;  wr_cycle[ 2316] = 1'b0;  addr_rom[ 2316]='h00000000;  wr_data_rom[ 2316]='h00000000;
    rd_cycle[ 2317] = 1'b0;  wr_cycle[ 2317] = 1'b0;  addr_rom[ 2317]='h00000000;  wr_data_rom[ 2317]='h00000000;
    rd_cycle[ 2318] = 1'b0;  wr_cycle[ 2318] = 1'b0;  addr_rom[ 2318]='h00000000;  wr_data_rom[ 2318]='h00000000;
    rd_cycle[ 2319] = 1'b0;  wr_cycle[ 2319] = 1'b0;  addr_rom[ 2319]='h00000000;  wr_data_rom[ 2319]='h00000000;
    rd_cycle[ 2320] = 1'b0;  wr_cycle[ 2320] = 1'b0;  addr_rom[ 2320]='h00000000;  wr_data_rom[ 2320]='h00000000;
    rd_cycle[ 2321] = 1'b0;  wr_cycle[ 2321] = 1'b0;  addr_rom[ 2321]='h00000000;  wr_data_rom[ 2321]='h00000000;
    rd_cycle[ 2322] = 1'b0;  wr_cycle[ 2322] = 1'b0;  addr_rom[ 2322]='h00000000;  wr_data_rom[ 2322]='h00000000;
    rd_cycle[ 2323] = 1'b0;  wr_cycle[ 2323] = 1'b0;  addr_rom[ 2323]='h00000000;  wr_data_rom[ 2323]='h00000000;
    rd_cycle[ 2324] = 1'b0;  wr_cycle[ 2324] = 1'b0;  addr_rom[ 2324]='h00000000;  wr_data_rom[ 2324]='h00000000;
    rd_cycle[ 2325] = 1'b0;  wr_cycle[ 2325] = 1'b0;  addr_rom[ 2325]='h00000000;  wr_data_rom[ 2325]='h00000000;
    rd_cycle[ 2326] = 1'b0;  wr_cycle[ 2326] = 1'b0;  addr_rom[ 2326]='h00000000;  wr_data_rom[ 2326]='h00000000;
    rd_cycle[ 2327] = 1'b0;  wr_cycle[ 2327] = 1'b0;  addr_rom[ 2327]='h00000000;  wr_data_rom[ 2327]='h00000000;
    rd_cycle[ 2328] = 1'b0;  wr_cycle[ 2328] = 1'b0;  addr_rom[ 2328]='h00000000;  wr_data_rom[ 2328]='h00000000;
    rd_cycle[ 2329] = 1'b0;  wr_cycle[ 2329] = 1'b0;  addr_rom[ 2329]='h00000000;  wr_data_rom[ 2329]='h00000000;
    rd_cycle[ 2330] = 1'b0;  wr_cycle[ 2330] = 1'b0;  addr_rom[ 2330]='h00000000;  wr_data_rom[ 2330]='h00000000;
    rd_cycle[ 2331] = 1'b0;  wr_cycle[ 2331] = 1'b0;  addr_rom[ 2331]='h00000000;  wr_data_rom[ 2331]='h00000000;
    rd_cycle[ 2332] = 1'b0;  wr_cycle[ 2332] = 1'b0;  addr_rom[ 2332]='h00000000;  wr_data_rom[ 2332]='h00000000;
    rd_cycle[ 2333] = 1'b0;  wr_cycle[ 2333] = 1'b0;  addr_rom[ 2333]='h00000000;  wr_data_rom[ 2333]='h00000000;
    rd_cycle[ 2334] = 1'b0;  wr_cycle[ 2334] = 1'b0;  addr_rom[ 2334]='h00000000;  wr_data_rom[ 2334]='h00000000;
    rd_cycle[ 2335] = 1'b0;  wr_cycle[ 2335] = 1'b0;  addr_rom[ 2335]='h00000000;  wr_data_rom[ 2335]='h00000000;
    rd_cycle[ 2336] = 1'b0;  wr_cycle[ 2336] = 1'b0;  addr_rom[ 2336]='h00000000;  wr_data_rom[ 2336]='h00000000;
    rd_cycle[ 2337] = 1'b0;  wr_cycle[ 2337] = 1'b0;  addr_rom[ 2337]='h00000000;  wr_data_rom[ 2337]='h00000000;
    rd_cycle[ 2338] = 1'b0;  wr_cycle[ 2338] = 1'b0;  addr_rom[ 2338]='h00000000;  wr_data_rom[ 2338]='h00000000;
    rd_cycle[ 2339] = 1'b0;  wr_cycle[ 2339] = 1'b0;  addr_rom[ 2339]='h00000000;  wr_data_rom[ 2339]='h00000000;
    rd_cycle[ 2340] = 1'b0;  wr_cycle[ 2340] = 1'b0;  addr_rom[ 2340]='h00000000;  wr_data_rom[ 2340]='h00000000;
    rd_cycle[ 2341] = 1'b0;  wr_cycle[ 2341] = 1'b0;  addr_rom[ 2341]='h00000000;  wr_data_rom[ 2341]='h00000000;
    rd_cycle[ 2342] = 1'b0;  wr_cycle[ 2342] = 1'b0;  addr_rom[ 2342]='h00000000;  wr_data_rom[ 2342]='h00000000;
    rd_cycle[ 2343] = 1'b0;  wr_cycle[ 2343] = 1'b0;  addr_rom[ 2343]='h00000000;  wr_data_rom[ 2343]='h00000000;
    rd_cycle[ 2344] = 1'b0;  wr_cycle[ 2344] = 1'b0;  addr_rom[ 2344]='h00000000;  wr_data_rom[ 2344]='h00000000;
    rd_cycle[ 2345] = 1'b0;  wr_cycle[ 2345] = 1'b0;  addr_rom[ 2345]='h00000000;  wr_data_rom[ 2345]='h00000000;
    rd_cycle[ 2346] = 1'b0;  wr_cycle[ 2346] = 1'b0;  addr_rom[ 2346]='h00000000;  wr_data_rom[ 2346]='h00000000;
    rd_cycle[ 2347] = 1'b0;  wr_cycle[ 2347] = 1'b0;  addr_rom[ 2347]='h00000000;  wr_data_rom[ 2347]='h00000000;
    rd_cycle[ 2348] = 1'b0;  wr_cycle[ 2348] = 1'b0;  addr_rom[ 2348]='h00000000;  wr_data_rom[ 2348]='h00000000;
    rd_cycle[ 2349] = 1'b0;  wr_cycle[ 2349] = 1'b0;  addr_rom[ 2349]='h00000000;  wr_data_rom[ 2349]='h00000000;
    rd_cycle[ 2350] = 1'b0;  wr_cycle[ 2350] = 1'b0;  addr_rom[ 2350]='h00000000;  wr_data_rom[ 2350]='h00000000;
    rd_cycle[ 2351] = 1'b0;  wr_cycle[ 2351] = 1'b0;  addr_rom[ 2351]='h00000000;  wr_data_rom[ 2351]='h00000000;
    rd_cycle[ 2352] = 1'b0;  wr_cycle[ 2352] = 1'b0;  addr_rom[ 2352]='h00000000;  wr_data_rom[ 2352]='h00000000;
    rd_cycle[ 2353] = 1'b0;  wr_cycle[ 2353] = 1'b0;  addr_rom[ 2353]='h00000000;  wr_data_rom[ 2353]='h00000000;
    rd_cycle[ 2354] = 1'b0;  wr_cycle[ 2354] = 1'b0;  addr_rom[ 2354]='h00000000;  wr_data_rom[ 2354]='h00000000;
    rd_cycle[ 2355] = 1'b0;  wr_cycle[ 2355] = 1'b0;  addr_rom[ 2355]='h00000000;  wr_data_rom[ 2355]='h00000000;
    rd_cycle[ 2356] = 1'b0;  wr_cycle[ 2356] = 1'b0;  addr_rom[ 2356]='h00000000;  wr_data_rom[ 2356]='h00000000;
    rd_cycle[ 2357] = 1'b0;  wr_cycle[ 2357] = 1'b0;  addr_rom[ 2357]='h00000000;  wr_data_rom[ 2357]='h00000000;
    rd_cycle[ 2358] = 1'b0;  wr_cycle[ 2358] = 1'b0;  addr_rom[ 2358]='h00000000;  wr_data_rom[ 2358]='h00000000;
    rd_cycle[ 2359] = 1'b0;  wr_cycle[ 2359] = 1'b0;  addr_rom[ 2359]='h00000000;  wr_data_rom[ 2359]='h00000000;
    rd_cycle[ 2360] = 1'b0;  wr_cycle[ 2360] = 1'b0;  addr_rom[ 2360]='h00000000;  wr_data_rom[ 2360]='h00000000;
    rd_cycle[ 2361] = 1'b0;  wr_cycle[ 2361] = 1'b0;  addr_rom[ 2361]='h00000000;  wr_data_rom[ 2361]='h00000000;
    rd_cycle[ 2362] = 1'b0;  wr_cycle[ 2362] = 1'b0;  addr_rom[ 2362]='h00000000;  wr_data_rom[ 2362]='h00000000;
    rd_cycle[ 2363] = 1'b0;  wr_cycle[ 2363] = 1'b0;  addr_rom[ 2363]='h00000000;  wr_data_rom[ 2363]='h00000000;
    rd_cycle[ 2364] = 1'b0;  wr_cycle[ 2364] = 1'b0;  addr_rom[ 2364]='h00000000;  wr_data_rom[ 2364]='h00000000;
    rd_cycle[ 2365] = 1'b0;  wr_cycle[ 2365] = 1'b0;  addr_rom[ 2365]='h00000000;  wr_data_rom[ 2365]='h00000000;
    rd_cycle[ 2366] = 1'b0;  wr_cycle[ 2366] = 1'b0;  addr_rom[ 2366]='h00000000;  wr_data_rom[ 2366]='h00000000;
    rd_cycle[ 2367] = 1'b0;  wr_cycle[ 2367] = 1'b0;  addr_rom[ 2367]='h00000000;  wr_data_rom[ 2367]='h00000000;
    rd_cycle[ 2368] = 1'b0;  wr_cycle[ 2368] = 1'b0;  addr_rom[ 2368]='h00000000;  wr_data_rom[ 2368]='h00000000;
    rd_cycle[ 2369] = 1'b0;  wr_cycle[ 2369] = 1'b0;  addr_rom[ 2369]='h00000000;  wr_data_rom[ 2369]='h00000000;
    rd_cycle[ 2370] = 1'b0;  wr_cycle[ 2370] = 1'b0;  addr_rom[ 2370]='h00000000;  wr_data_rom[ 2370]='h00000000;
    rd_cycle[ 2371] = 1'b0;  wr_cycle[ 2371] = 1'b0;  addr_rom[ 2371]='h00000000;  wr_data_rom[ 2371]='h00000000;
    rd_cycle[ 2372] = 1'b0;  wr_cycle[ 2372] = 1'b0;  addr_rom[ 2372]='h00000000;  wr_data_rom[ 2372]='h00000000;
    rd_cycle[ 2373] = 1'b0;  wr_cycle[ 2373] = 1'b0;  addr_rom[ 2373]='h00000000;  wr_data_rom[ 2373]='h00000000;
    rd_cycle[ 2374] = 1'b0;  wr_cycle[ 2374] = 1'b0;  addr_rom[ 2374]='h00000000;  wr_data_rom[ 2374]='h00000000;
    rd_cycle[ 2375] = 1'b0;  wr_cycle[ 2375] = 1'b0;  addr_rom[ 2375]='h00000000;  wr_data_rom[ 2375]='h00000000;
    rd_cycle[ 2376] = 1'b0;  wr_cycle[ 2376] = 1'b0;  addr_rom[ 2376]='h00000000;  wr_data_rom[ 2376]='h00000000;
    rd_cycle[ 2377] = 1'b0;  wr_cycle[ 2377] = 1'b0;  addr_rom[ 2377]='h00000000;  wr_data_rom[ 2377]='h00000000;
    rd_cycle[ 2378] = 1'b0;  wr_cycle[ 2378] = 1'b0;  addr_rom[ 2378]='h00000000;  wr_data_rom[ 2378]='h00000000;
    rd_cycle[ 2379] = 1'b0;  wr_cycle[ 2379] = 1'b0;  addr_rom[ 2379]='h00000000;  wr_data_rom[ 2379]='h00000000;
    rd_cycle[ 2380] = 1'b0;  wr_cycle[ 2380] = 1'b0;  addr_rom[ 2380]='h00000000;  wr_data_rom[ 2380]='h00000000;
    rd_cycle[ 2381] = 1'b0;  wr_cycle[ 2381] = 1'b0;  addr_rom[ 2381]='h00000000;  wr_data_rom[ 2381]='h00000000;
    rd_cycle[ 2382] = 1'b0;  wr_cycle[ 2382] = 1'b0;  addr_rom[ 2382]='h00000000;  wr_data_rom[ 2382]='h00000000;
    rd_cycle[ 2383] = 1'b0;  wr_cycle[ 2383] = 1'b0;  addr_rom[ 2383]='h00000000;  wr_data_rom[ 2383]='h00000000;
    rd_cycle[ 2384] = 1'b0;  wr_cycle[ 2384] = 1'b0;  addr_rom[ 2384]='h00000000;  wr_data_rom[ 2384]='h00000000;
    rd_cycle[ 2385] = 1'b0;  wr_cycle[ 2385] = 1'b0;  addr_rom[ 2385]='h00000000;  wr_data_rom[ 2385]='h00000000;
    rd_cycle[ 2386] = 1'b0;  wr_cycle[ 2386] = 1'b0;  addr_rom[ 2386]='h00000000;  wr_data_rom[ 2386]='h00000000;
    rd_cycle[ 2387] = 1'b0;  wr_cycle[ 2387] = 1'b0;  addr_rom[ 2387]='h00000000;  wr_data_rom[ 2387]='h00000000;
    rd_cycle[ 2388] = 1'b0;  wr_cycle[ 2388] = 1'b0;  addr_rom[ 2388]='h00000000;  wr_data_rom[ 2388]='h00000000;
    rd_cycle[ 2389] = 1'b0;  wr_cycle[ 2389] = 1'b0;  addr_rom[ 2389]='h00000000;  wr_data_rom[ 2389]='h00000000;
    rd_cycle[ 2390] = 1'b0;  wr_cycle[ 2390] = 1'b0;  addr_rom[ 2390]='h00000000;  wr_data_rom[ 2390]='h00000000;
    rd_cycle[ 2391] = 1'b0;  wr_cycle[ 2391] = 1'b0;  addr_rom[ 2391]='h00000000;  wr_data_rom[ 2391]='h00000000;
    rd_cycle[ 2392] = 1'b0;  wr_cycle[ 2392] = 1'b0;  addr_rom[ 2392]='h00000000;  wr_data_rom[ 2392]='h00000000;
    rd_cycle[ 2393] = 1'b0;  wr_cycle[ 2393] = 1'b0;  addr_rom[ 2393]='h00000000;  wr_data_rom[ 2393]='h00000000;
    rd_cycle[ 2394] = 1'b0;  wr_cycle[ 2394] = 1'b0;  addr_rom[ 2394]='h00000000;  wr_data_rom[ 2394]='h00000000;
    rd_cycle[ 2395] = 1'b0;  wr_cycle[ 2395] = 1'b0;  addr_rom[ 2395]='h00000000;  wr_data_rom[ 2395]='h00000000;
    rd_cycle[ 2396] = 1'b0;  wr_cycle[ 2396] = 1'b0;  addr_rom[ 2396]='h00000000;  wr_data_rom[ 2396]='h00000000;
    rd_cycle[ 2397] = 1'b0;  wr_cycle[ 2397] = 1'b0;  addr_rom[ 2397]='h00000000;  wr_data_rom[ 2397]='h00000000;
    rd_cycle[ 2398] = 1'b0;  wr_cycle[ 2398] = 1'b0;  addr_rom[ 2398]='h00000000;  wr_data_rom[ 2398]='h00000000;
    rd_cycle[ 2399] = 1'b0;  wr_cycle[ 2399] = 1'b0;  addr_rom[ 2399]='h00000000;  wr_data_rom[ 2399]='h00000000;
    rd_cycle[ 2400] = 1'b0;  wr_cycle[ 2400] = 1'b0;  addr_rom[ 2400]='h00000000;  wr_data_rom[ 2400]='h00000000;
    rd_cycle[ 2401] = 1'b0;  wr_cycle[ 2401] = 1'b0;  addr_rom[ 2401]='h00000000;  wr_data_rom[ 2401]='h00000000;
    rd_cycle[ 2402] = 1'b0;  wr_cycle[ 2402] = 1'b0;  addr_rom[ 2402]='h00000000;  wr_data_rom[ 2402]='h00000000;
    rd_cycle[ 2403] = 1'b0;  wr_cycle[ 2403] = 1'b0;  addr_rom[ 2403]='h00000000;  wr_data_rom[ 2403]='h00000000;
    rd_cycle[ 2404] = 1'b0;  wr_cycle[ 2404] = 1'b0;  addr_rom[ 2404]='h00000000;  wr_data_rom[ 2404]='h00000000;
    rd_cycle[ 2405] = 1'b0;  wr_cycle[ 2405] = 1'b0;  addr_rom[ 2405]='h00000000;  wr_data_rom[ 2405]='h00000000;
    rd_cycle[ 2406] = 1'b0;  wr_cycle[ 2406] = 1'b0;  addr_rom[ 2406]='h00000000;  wr_data_rom[ 2406]='h00000000;
    rd_cycle[ 2407] = 1'b0;  wr_cycle[ 2407] = 1'b0;  addr_rom[ 2407]='h00000000;  wr_data_rom[ 2407]='h00000000;
    rd_cycle[ 2408] = 1'b0;  wr_cycle[ 2408] = 1'b0;  addr_rom[ 2408]='h00000000;  wr_data_rom[ 2408]='h00000000;
    rd_cycle[ 2409] = 1'b0;  wr_cycle[ 2409] = 1'b0;  addr_rom[ 2409]='h00000000;  wr_data_rom[ 2409]='h00000000;
    rd_cycle[ 2410] = 1'b0;  wr_cycle[ 2410] = 1'b0;  addr_rom[ 2410]='h00000000;  wr_data_rom[ 2410]='h00000000;
    rd_cycle[ 2411] = 1'b0;  wr_cycle[ 2411] = 1'b0;  addr_rom[ 2411]='h00000000;  wr_data_rom[ 2411]='h00000000;
    rd_cycle[ 2412] = 1'b0;  wr_cycle[ 2412] = 1'b0;  addr_rom[ 2412]='h00000000;  wr_data_rom[ 2412]='h00000000;
    rd_cycle[ 2413] = 1'b0;  wr_cycle[ 2413] = 1'b0;  addr_rom[ 2413]='h00000000;  wr_data_rom[ 2413]='h00000000;
    rd_cycle[ 2414] = 1'b0;  wr_cycle[ 2414] = 1'b0;  addr_rom[ 2414]='h00000000;  wr_data_rom[ 2414]='h00000000;
    rd_cycle[ 2415] = 1'b0;  wr_cycle[ 2415] = 1'b0;  addr_rom[ 2415]='h00000000;  wr_data_rom[ 2415]='h00000000;
    rd_cycle[ 2416] = 1'b0;  wr_cycle[ 2416] = 1'b0;  addr_rom[ 2416]='h00000000;  wr_data_rom[ 2416]='h00000000;
    rd_cycle[ 2417] = 1'b0;  wr_cycle[ 2417] = 1'b0;  addr_rom[ 2417]='h00000000;  wr_data_rom[ 2417]='h00000000;
    rd_cycle[ 2418] = 1'b0;  wr_cycle[ 2418] = 1'b0;  addr_rom[ 2418]='h00000000;  wr_data_rom[ 2418]='h00000000;
    rd_cycle[ 2419] = 1'b0;  wr_cycle[ 2419] = 1'b0;  addr_rom[ 2419]='h00000000;  wr_data_rom[ 2419]='h00000000;
    rd_cycle[ 2420] = 1'b0;  wr_cycle[ 2420] = 1'b0;  addr_rom[ 2420]='h00000000;  wr_data_rom[ 2420]='h00000000;
    rd_cycle[ 2421] = 1'b0;  wr_cycle[ 2421] = 1'b0;  addr_rom[ 2421]='h00000000;  wr_data_rom[ 2421]='h00000000;
    rd_cycle[ 2422] = 1'b0;  wr_cycle[ 2422] = 1'b0;  addr_rom[ 2422]='h00000000;  wr_data_rom[ 2422]='h00000000;
    rd_cycle[ 2423] = 1'b0;  wr_cycle[ 2423] = 1'b0;  addr_rom[ 2423]='h00000000;  wr_data_rom[ 2423]='h00000000;
    rd_cycle[ 2424] = 1'b0;  wr_cycle[ 2424] = 1'b0;  addr_rom[ 2424]='h00000000;  wr_data_rom[ 2424]='h00000000;
    rd_cycle[ 2425] = 1'b0;  wr_cycle[ 2425] = 1'b0;  addr_rom[ 2425]='h00000000;  wr_data_rom[ 2425]='h00000000;
    rd_cycle[ 2426] = 1'b0;  wr_cycle[ 2426] = 1'b0;  addr_rom[ 2426]='h00000000;  wr_data_rom[ 2426]='h00000000;
    rd_cycle[ 2427] = 1'b0;  wr_cycle[ 2427] = 1'b0;  addr_rom[ 2427]='h00000000;  wr_data_rom[ 2427]='h00000000;
    rd_cycle[ 2428] = 1'b0;  wr_cycle[ 2428] = 1'b0;  addr_rom[ 2428]='h00000000;  wr_data_rom[ 2428]='h00000000;
    rd_cycle[ 2429] = 1'b0;  wr_cycle[ 2429] = 1'b0;  addr_rom[ 2429]='h00000000;  wr_data_rom[ 2429]='h00000000;
    rd_cycle[ 2430] = 1'b0;  wr_cycle[ 2430] = 1'b0;  addr_rom[ 2430]='h00000000;  wr_data_rom[ 2430]='h00000000;
    rd_cycle[ 2431] = 1'b0;  wr_cycle[ 2431] = 1'b0;  addr_rom[ 2431]='h00000000;  wr_data_rom[ 2431]='h00000000;
    rd_cycle[ 2432] = 1'b0;  wr_cycle[ 2432] = 1'b0;  addr_rom[ 2432]='h00000000;  wr_data_rom[ 2432]='h00000000;
    rd_cycle[ 2433] = 1'b0;  wr_cycle[ 2433] = 1'b0;  addr_rom[ 2433]='h00000000;  wr_data_rom[ 2433]='h00000000;
    rd_cycle[ 2434] = 1'b0;  wr_cycle[ 2434] = 1'b0;  addr_rom[ 2434]='h00000000;  wr_data_rom[ 2434]='h00000000;
    rd_cycle[ 2435] = 1'b0;  wr_cycle[ 2435] = 1'b0;  addr_rom[ 2435]='h00000000;  wr_data_rom[ 2435]='h00000000;
    rd_cycle[ 2436] = 1'b0;  wr_cycle[ 2436] = 1'b0;  addr_rom[ 2436]='h00000000;  wr_data_rom[ 2436]='h00000000;
    rd_cycle[ 2437] = 1'b0;  wr_cycle[ 2437] = 1'b0;  addr_rom[ 2437]='h00000000;  wr_data_rom[ 2437]='h00000000;
    rd_cycle[ 2438] = 1'b0;  wr_cycle[ 2438] = 1'b0;  addr_rom[ 2438]='h00000000;  wr_data_rom[ 2438]='h00000000;
    rd_cycle[ 2439] = 1'b0;  wr_cycle[ 2439] = 1'b0;  addr_rom[ 2439]='h00000000;  wr_data_rom[ 2439]='h00000000;
    rd_cycle[ 2440] = 1'b0;  wr_cycle[ 2440] = 1'b0;  addr_rom[ 2440]='h00000000;  wr_data_rom[ 2440]='h00000000;
    rd_cycle[ 2441] = 1'b0;  wr_cycle[ 2441] = 1'b0;  addr_rom[ 2441]='h00000000;  wr_data_rom[ 2441]='h00000000;
    rd_cycle[ 2442] = 1'b0;  wr_cycle[ 2442] = 1'b0;  addr_rom[ 2442]='h00000000;  wr_data_rom[ 2442]='h00000000;
    rd_cycle[ 2443] = 1'b0;  wr_cycle[ 2443] = 1'b0;  addr_rom[ 2443]='h00000000;  wr_data_rom[ 2443]='h00000000;
    rd_cycle[ 2444] = 1'b0;  wr_cycle[ 2444] = 1'b0;  addr_rom[ 2444]='h00000000;  wr_data_rom[ 2444]='h00000000;
    rd_cycle[ 2445] = 1'b0;  wr_cycle[ 2445] = 1'b0;  addr_rom[ 2445]='h00000000;  wr_data_rom[ 2445]='h00000000;
    rd_cycle[ 2446] = 1'b0;  wr_cycle[ 2446] = 1'b0;  addr_rom[ 2446]='h00000000;  wr_data_rom[ 2446]='h00000000;
    rd_cycle[ 2447] = 1'b0;  wr_cycle[ 2447] = 1'b0;  addr_rom[ 2447]='h00000000;  wr_data_rom[ 2447]='h00000000;
    rd_cycle[ 2448] = 1'b0;  wr_cycle[ 2448] = 1'b0;  addr_rom[ 2448]='h00000000;  wr_data_rom[ 2448]='h00000000;
    rd_cycle[ 2449] = 1'b0;  wr_cycle[ 2449] = 1'b0;  addr_rom[ 2449]='h00000000;  wr_data_rom[ 2449]='h00000000;
    rd_cycle[ 2450] = 1'b0;  wr_cycle[ 2450] = 1'b0;  addr_rom[ 2450]='h00000000;  wr_data_rom[ 2450]='h00000000;
    rd_cycle[ 2451] = 1'b0;  wr_cycle[ 2451] = 1'b0;  addr_rom[ 2451]='h00000000;  wr_data_rom[ 2451]='h00000000;
    rd_cycle[ 2452] = 1'b0;  wr_cycle[ 2452] = 1'b0;  addr_rom[ 2452]='h00000000;  wr_data_rom[ 2452]='h00000000;
    rd_cycle[ 2453] = 1'b0;  wr_cycle[ 2453] = 1'b0;  addr_rom[ 2453]='h00000000;  wr_data_rom[ 2453]='h00000000;
    rd_cycle[ 2454] = 1'b0;  wr_cycle[ 2454] = 1'b0;  addr_rom[ 2454]='h00000000;  wr_data_rom[ 2454]='h00000000;
    rd_cycle[ 2455] = 1'b0;  wr_cycle[ 2455] = 1'b0;  addr_rom[ 2455]='h00000000;  wr_data_rom[ 2455]='h00000000;
    rd_cycle[ 2456] = 1'b0;  wr_cycle[ 2456] = 1'b0;  addr_rom[ 2456]='h00000000;  wr_data_rom[ 2456]='h00000000;
    rd_cycle[ 2457] = 1'b0;  wr_cycle[ 2457] = 1'b0;  addr_rom[ 2457]='h00000000;  wr_data_rom[ 2457]='h00000000;
    rd_cycle[ 2458] = 1'b0;  wr_cycle[ 2458] = 1'b0;  addr_rom[ 2458]='h00000000;  wr_data_rom[ 2458]='h00000000;
    rd_cycle[ 2459] = 1'b0;  wr_cycle[ 2459] = 1'b0;  addr_rom[ 2459]='h00000000;  wr_data_rom[ 2459]='h00000000;
    rd_cycle[ 2460] = 1'b0;  wr_cycle[ 2460] = 1'b0;  addr_rom[ 2460]='h00000000;  wr_data_rom[ 2460]='h00000000;
    rd_cycle[ 2461] = 1'b0;  wr_cycle[ 2461] = 1'b0;  addr_rom[ 2461]='h00000000;  wr_data_rom[ 2461]='h00000000;
    rd_cycle[ 2462] = 1'b0;  wr_cycle[ 2462] = 1'b0;  addr_rom[ 2462]='h00000000;  wr_data_rom[ 2462]='h00000000;
    rd_cycle[ 2463] = 1'b0;  wr_cycle[ 2463] = 1'b0;  addr_rom[ 2463]='h00000000;  wr_data_rom[ 2463]='h00000000;
    rd_cycle[ 2464] = 1'b0;  wr_cycle[ 2464] = 1'b0;  addr_rom[ 2464]='h00000000;  wr_data_rom[ 2464]='h00000000;
    rd_cycle[ 2465] = 1'b0;  wr_cycle[ 2465] = 1'b0;  addr_rom[ 2465]='h00000000;  wr_data_rom[ 2465]='h00000000;
    rd_cycle[ 2466] = 1'b0;  wr_cycle[ 2466] = 1'b0;  addr_rom[ 2466]='h00000000;  wr_data_rom[ 2466]='h00000000;
    rd_cycle[ 2467] = 1'b0;  wr_cycle[ 2467] = 1'b0;  addr_rom[ 2467]='h00000000;  wr_data_rom[ 2467]='h00000000;
    rd_cycle[ 2468] = 1'b0;  wr_cycle[ 2468] = 1'b0;  addr_rom[ 2468]='h00000000;  wr_data_rom[ 2468]='h00000000;
    rd_cycle[ 2469] = 1'b0;  wr_cycle[ 2469] = 1'b0;  addr_rom[ 2469]='h00000000;  wr_data_rom[ 2469]='h00000000;
    rd_cycle[ 2470] = 1'b0;  wr_cycle[ 2470] = 1'b0;  addr_rom[ 2470]='h00000000;  wr_data_rom[ 2470]='h00000000;
    rd_cycle[ 2471] = 1'b0;  wr_cycle[ 2471] = 1'b0;  addr_rom[ 2471]='h00000000;  wr_data_rom[ 2471]='h00000000;
    rd_cycle[ 2472] = 1'b0;  wr_cycle[ 2472] = 1'b0;  addr_rom[ 2472]='h00000000;  wr_data_rom[ 2472]='h00000000;
    rd_cycle[ 2473] = 1'b0;  wr_cycle[ 2473] = 1'b0;  addr_rom[ 2473]='h00000000;  wr_data_rom[ 2473]='h00000000;
    rd_cycle[ 2474] = 1'b0;  wr_cycle[ 2474] = 1'b0;  addr_rom[ 2474]='h00000000;  wr_data_rom[ 2474]='h00000000;
    rd_cycle[ 2475] = 1'b0;  wr_cycle[ 2475] = 1'b0;  addr_rom[ 2475]='h00000000;  wr_data_rom[ 2475]='h00000000;
    rd_cycle[ 2476] = 1'b0;  wr_cycle[ 2476] = 1'b0;  addr_rom[ 2476]='h00000000;  wr_data_rom[ 2476]='h00000000;
    rd_cycle[ 2477] = 1'b0;  wr_cycle[ 2477] = 1'b0;  addr_rom[ 2477]='h00000000;  wr_data_rom[ 2477]='h00000000;
    rd_cycle[ 2478] = 1'b0;  wr_cycle[ 2478] = 1'b0;  addr_rom[ 2478]='h00000000;  wr_data_rom[ 2478]='h00000000;
    rd_cycle[ 2479] = 1'b0;  wr_cycle[ 2479] = 1'b0;  addr_rom[ 2479]='h00000000;  wr_data_rom[ 2479]='h00000000;
    rd_cycle[ 2480] = 1'b0;  wr_cycle[ 2480] = 1'b0;  addr_rom[ 2480]='h00000000;  wr_data_rom[ 2480]='h00000000;
    rd_cycle[ 2481] = 1'b0;  wr_cycle[ 2481] = 1'b0;  addr_rom[ 2481]='h00000000;  wr_data_rom[ 2481]='h00000000;
    rd_cycle[ 2482] = 1'b0;  wr_cycle[ 2482] = 1'b0;  addr_rom[ 2482]='h00000000;  wr_data_rom[ 2482]='h00000000;
    rd_cycle[ 2483] = 1'b0;  wr_cycle[ 2483] = 1'b0;  addr_rom[ 2483]='h00000000;  wr_data_rom[ 2483]='h00000000;
    rd_cycle[ 2484] = 1'b0;  wr_cycle[ 2484] = 1'b0;  addr_rom[ 2484]='h00000000;  wr_data_rom[ 2484]='h00000000;
    rd_cycle[ 2485] = 1'b0;  wr_cycle[ 2485] = 1'b0;  addr_rom[ 2485]='h00000000;  wr_data_rom[ 2485]='h00000000;
    rd_cycle[ 2486] = 1'b0;  wr_cycle[ 2486] = 1'b0;  addr_rom[ 2486]='h00000000;  wr_data_rom[ 2486]='h00000000;
    rd_cycle[ 2487] = 1'b0;  wr_cycle[ 2487] = 1'b0;  addr_rom[ 2487]='h00000000;  wr_data_rom[ 2487]='h00000000;
    rd_cycle[ 2488] = 1'b0;  wr_cycle[ 2488] = 1'b0;  addr_rom[ 2488]='h00000000;  wr_data_rom[ 2488]='h00000000;
    rd_cycle[ 2489] = 1'b0;  wr_cycle[ 2489] = 1'b0;  addr_rom[ 2489]='h00000000;  wr_data_rom[ 2489]='h00000000;
    rd_cycle[ 2490] = 1'b0;  wr_cycle[ 2490] = 1'b0;  addr_rom[ 2490]='h00000000;  wr_data_rom[ 2490]='h00000000;
    rd_cycle[ 2491] = 1'b0;  wr_cycle[ 2491] = 1'b0;  addr_rom[ 2491]='h00000000;  wr_data_rom[ 2491]='h00000000;
    rd_cycle[ 2492] = 1'b0;  wr_cycle[ 2492] = 1'b0;  addr_rom[ 2492]='h00000000;  wr_data_rom[ 2492]='h00000000;
    rd_cycle[ 2493] = 1'b0;  wr_cycle[ 2493] = 1'b0;  addr_rom[ 2493]='h00000000;  wr_data_rom[ 2493]='h00000000;
    rd_cycle[ 2494] = 1'b0;  wr_cycle[ 2494] = 1'b0;  addr_rom[ 2494]='h00000000;  wr_data_rom[ 2494]='h00000000;
    rd_cycle[ 2495] = 1'b0;  wr_cycle[ 2495] = 1'b0;  addr_rom[ 2495]='h00000000;  wr_data_rom[ 2495]='h00000000;
    rd_cycle[ 2496] = 1'b0;  wr_cycle[ 2496] = 1'b0;  addr_rom[ 2496]='h00000000;  wr_data_rom[ 2496]='h00000000;
    rd_cycle[ 2497] = 1'b0;  wr_cycle[ 2497] = 1'b0;  addr_rom[ 2497]='h00000000;  wr_data_rom[ 2497]='h00000000;
    rd_cycle[ 2498] = 1'b0;  wr_cycle[ 2498] = 1'b0;  addr_rom[ 2498]='h00000000;  wr_data_rom[ 2498]='h00000000;
    rd_cycle[ 2499] = 1'b0;  wr_cycle[ 2499] = 1'b0;  addr_rom[ 2499]='h00000000;  wr_data_rom[ 2499]='h00000000;
    rd_cycle[ 2500] = 1'b0;  wr_cycle[ 2500] = 1'b0;  addr_rom[ 2500]='h00000000;  wr_data_rom[ 2500]='h00000000;
    rd_cycle[ 2501] = 1'b0;  wr_cycle[ 2501] = 1'b0;  addr_rom[ 2501]='h00000000;  wr_data_rom[ 2501]='h00000000;
    rd_cycle[ 2502] = 1'b0;  wr_cycle[ 2502] = 1'b0;  addr_rom[ 2502]='h00000000;  wr_data_rom[ 2502]='h00000000;
    rd_cycle[ 2503] = 1'b0;  wr_cycle[ 2503] = 1'b0;  addr_rom[ 2503]='h00000000;  wr_data_rom[ 2503]='h00000000;
    rd_cycle[ 2504] = 1'b0;  wr_cycle[ 2504] = 1'b0;  addr_rom[ 2504]='h00000000;  wr_data_rom[ 2504]='h00000000;
    rd_cycle[ 2505] = 1'b0;  wr_cycle[ 2505] = 1'b0;  addr_rom[ 2505]='h00000000;  wr_data_rom[ 2505]='h00000000;
    rd_cycle[ 2506] = 1'b0;  wr_cycle[ 2506] = 1'b0;  addr_rom[ 2506]='h00000000;  wr_data_rom[ 2506]='h00000000;
    rd_cycle[ 2507] = 1'b0;  wr_cycle[ 2507] = 1'b0;  addr_rom[ 2507]='h00000000;  wr_data_rom[ 2507]='h00000000;
    rd_cycle[ 2508] = 1'b0;  wr_cycle[ 2508] = 1'b0;  addr_rom[ 2508]='h00000000;  wr_data_rom[ 2508]='h00000000;
    rd_cycle[ 2509] = 1'b0;  wr_cycle[ 2509] = 1'b0;  addr_rom[ 2509]='h00000000;  wr_data_rom[ 2509]='h00000000;
    rd_cycle[ 2510] = 1'b0;  wr_cycle[ 2510] = 1'b0;  addr_rom[ 2510]='h00000000;  wr_data_rom[ 2510]='h00000000;
    rd_cycle[ 2511] = 1'b0;  wr_cycle[ 2511] = 1'b0;  addr_rom[ 2511]='h00000000;  wr_data_rom[ 2511]='h00000000;
    rd_cycle[ 2512] = 1'b0;  wr_cycle[ 2512] = 1'b0;  addr_rom[ 2512]='h00000000;  wr_data_rom[ 2512]='h00000000;
    rd_cycle[ 2513] = 1'b0;  wr_cycle[ 2513] = 1'b0;  addr_rom[ 2513]='h00000000;  wr_data_rom[ 2513]='h00000000;
    rd_cycle[ 2514] = 1'b0;  wr_cycle[ 2514] = 1'b0;  addr_rom[ 2514]='h00000000;  wr_data_rom[ 2514]='h00000000;
    rd_cycle[ 2515] = 1'b0;  wr_cycle[ 2515] = 1'b0;  addr_rom[ 2515]='h00000000;  wr_data_rom[ 2515]='h00000000;
    rd_cycle[ 2516] = 1'b0;  wr_cycle[ 2516] = 1'b0;  addr_rom[ 2516]='h00000000;  wr_data_rom[ 2516]='h00000000;
    rd_cycle[ 2517] = 1'b0;  wr_cycle[ 2517] = 1'b0;  addr_rom[ 2517]='h00000000;  wr_data_rom[ 2517]='h00000000;
    rd_cycle[ 2518] = 1'b0;  wr_cycle[ 2518] = 1'b0;  addr_rom[ 2518]='h00000000;  wr_data_rom[ 2518]='h00000000;
    rd_cycle[ 2519] = 1'b0;  wr_cycle[ 2519] = 1'b0;  addr_rom[ 2519]='h00000000;  wr_data_rom[ 2519]='h00000000;
    rd_cycle[ 2520] = 1'b0;  wr_cycle[ 2520] = 1'b0;  addr_rom[ 2520]='h00000000;  wr_data_rom[ 2520]='h00000000;
    rd_cycle[ 2521] = 1'b0;  wr_cycle[ 2521] = 1'b0;  addr_rom[ 2521]='h00000000;  wr_data_rom[ 2521]='h00000000;
    rd_cycle[ 2522] = 1'b0;  wr_cycle[ 2522] = 1'b0;  addr_rom[ 2522]='h00000000;  wr_data_rom[ 2522]='h00000000;
    rd_cycle[ 2523] = 1'b0;  wr_cycle[ 2523] = 1'b0;  addr_rom[ 2523]='h00000000;  wr_data_rom[ 2523]='h00000000;
    rd_cycle[ 2524] = 1'b0;  wr_cycle[ 2524] = 1'b0;  addr_rom[ 2524]='h00000000;  wr_data_rom[ 2524]='h00000000;
    rd_cycle[ 2525] = 1'b0;  wr_cycle[ 2525] = 1'b0;  addr_rom[ 2525]='h00000000;  wr_data_rom[ 2525]='h00000000;
    rd_cycle[ 2526] = 1'b0;  wr_cycle[ 2526] = 1'b0;  addr_rom[ 2526]='h00000000;  wr_data_rom[ 2526]='h00000000;
    rd_cycle[ 2527] = 1'b0;  wr_cycle[ 2527] = 1'b0;  addr_rom[ 2527]='h00000000;  wr_data_rom[ 2527]='h00000000;
    rd_cycle[ 2528] = 1'b0;  wr_cycle[ 2528] = 1'b0;  addr_rom[ 2528]='h00000000;  wr_data_rom[ 2528]='h00000000;
    rd_cycle[ 2529] = 1'b0;  wr_cycle[ 2529] = 1'b0;  addr_rom[ 2529]='h00000000;  wr_data_rom[ 2529]='h00000000;
    rd_cycle[ 2530] = 1'b0;  wr_cycle[ 2530] = 1'b0;  addr_rom[ 2530]='h00000000;  wr_data_rom[ 2530]='h00000000;
    rd_cycle[ 2531] = 1'b0;  wr_cycle[ 2531] = 1'b0;  addr_rom[ 2531]='h00000000;  wr_data_rom[ 2531]='h00000000;
    rd_cycle[ 2532] = 1'b0;  wr_cycle[ 2532] = 1'b0;  addr_rom[ 2532]='h00000000;  wr_data_rom[ 2532]='h00000000;
    rd_cycle[ 2533] = 1'b0;  wr_cycle[ 2533] = 1'b0;  addr_rom[ 2533]='h00000000;  wr_data_rom[ 2533]='h00000000;
    rd_cycle[ 2534] = 1'b0;  wr_cycle[ 2534] = 1'b0;  addr_rom[ 2534]='h00000000;  wr_data_rom[ 2534]='h00000000;
    rd_cycle[ 2535] = 1'b0;  wr_cycle[ 2535] = 1'b0;  addr_rom[ 2535]='h00000000;  wr_data_rom[ 2535]='h00000000;
    rd_cycle[ 2536] = 1'b0;  wr_cycle[ 2536] = 1'b0;  addr_rom[ 2536]='h00000000;  wr_data_rom[ 2536]='h00000000;
    rd_cycle[ 2537] = 1'b0;  wr_cycle[ 2537] = 1'b0;  addr_rom[ 2537]='h00000000;  wr_data_rom[ 2537]='h00000000;
    rd_cycle[ 2538] = 1'b0;  wr_cycle[ 2538] = 1'b0;  addr_rom[ 2538]='h00000000;  wr_data_rom[ 2538]='h00000000;
    rd_cycle[ 2539] = 1'b0;  wr_cycle[ 2539] = 1'b0;  addr_rom[ 2539]='h00000000;  wr_data_rom[ 2539]='h00000000;
    rd_cycle[ 2540] = 1'b0;  wr_cycle[ 2540] = 1'b0;  addr_rom[ 2540]='h00000000;  wr_data_rom[ 2540]='h00000000;
    rd_cycle[ 2541] = 1'b0;  wr_cycle[ 2541] = 1'b0;  addr_rom[ 2541]='h00000000;  wr_data_rom[ 2541]='h00000000;
    rd_cycle[ 2542] = 1'b0;  wr_cycle[ 2542] = 1'b0;  addr_rom[ 2542]='h00000000;  wr_data_rom[ 2542]='h00000000;
    rd_cycle[ 2543] = 1'b0;  wr_cycle[ 2543] = 1'b0;  addr_rom[ 2543]='h00000000;  wr_data_rom[ 2543]='h00000000;
    rd_cycle[ 2544] = 1'b0;  wr_cycle[ 2544] = 1'b0;  addr_rom[ 2544]='h00000000;  wr_data_rom[ 2544]='h00000000;
    rd_cycle[ 2545] = 1'b0;  wr_cycle[ 2545] = 1'b0;  addr_rom[ 2545]='h00000000;  wr_data_rom[ 2545]='h00000000;
    rd_cycle[ 2546] = 1'b0;  wr_cycle[ 2546] = 1'b0;  addr_rom[ 2546]='h00000000;  wr_data_rom[ 2546]='h00000000;
    rd_cycle[ 2547] = 1'b0;  wr_cycle[ 2547] = 1'b0;  addr_rom[ 2547]='h00000000;  wr_data_rom[ 2547]='h00000000;
    rd_cycle[ 2548] = 1'b0;  wr_cycle[ 2548] = 1'b0;  addr_rom[ 2548]='h00000000;  wr_data_rom[ 2548]='h00000000;
    rd_cycle[ 2549] = 1'b0;  wr_cycle[ 2549] = 1'b0;  addr_rom[ 2549]='h00000000;  wr_data_rom[ 2549]='h00000000;
    rd_cycle[ 2550] = 1'b0;  wr_cycle[ 2550] = 1'b0;  addr_rom[ 2550]='h00000000;  wr_data_rom[ 2550]='h00000000;
    rd_cycle[ 2551] = 1'b0;  wr_cycle[ 2551] = 1'b0;  addr_rom[ 2551]='h00000000;  wr_data_rom[ 2551]='h00000000;
    rd_cycle[ 2552] = 1'b0;  wr_cycle[ 2552] = 1'b0;  addr_rom[ 2552]='h00000000;  wr_data_rom[ 2552]='h00000000;
    rd_cycle[ 2553] = 1'b0;  wr_cycle[ 2553] = 1'b0;  addr_rom[ 2553]='h00000000;  wr_data_rom[ 2553]='h00000000;
    rd_cycle[ 2554] = 1'b0;  wr_cycle[ 2554] = 1'b0;  addr_rom[ 2554]='h00000000;  wr_data_rom[ 2554]='h00000000;
    rd_cycle[ 2555] = 1'b0;  wr_cycle[ 2555] = 1'b0;  addr_rom[ 2555]='h00000000;  wr_data_rom[ 2555]='h00000000;
    rd_cycle[ 2556] = 1'b0;  wr_cycle[ 2556] = 1'b0;  addr_rom[ 2556]='h00000000;  wr_data_rom[ 2556]='h00000000;
    rd_cycle[ 2557] = 1'b0;  wr_cycle[ 2557] = 1'b0;  addr_rom[ 2557]='h00000000;  wr_data_rom[ 2557]='h00000000;
    rd_cycle[ 2558] = 1'b0;  wr_cycle[ 2558] = 1'b0;  addr_rom[ 2558]='h00000000;  wr_data_rom[ 2558]='h00000000;
    rd_cycle[ 2559] = 1'b0;  wr_cycle[ 2559] = 1'b0;  addr_rom[ 2559]='h00000000;  wr_data_rom[ 2559]='h00000000;
    // 512 sequence read cycles
    rd_cycle[ 2560] = 1'b1;  wr_cycle[ 2560] = 1'b0;  addr_rom[ 2560]='h00000000;  wr_data_rom[ 2560]='h00000000;
    rd_cycle[ 2561] = 1'b1;  wr_cycle[ 2561] = 1'b0;  addr_rom[ 2561]='h00000004;  wr_data_rom[ 2561]='h00000000;
    rd_cycle[ 2562] = 1'b1;  wr_cycle[ 2562] = 1'b0;  addr_rom[ 2562]='h00000008;  wr_data_rom[ 2562]='h00000000;
    rd_cycle[ 2563] = 1'b1;  wr_cycle[ 2563] = 1'b0;  addr_rom[ 2563]='h0000000c;  wr_data_rom[ 2563]='h00000000;
    rd_cycle[ 2564] = 1'b1;  wr_cycle[ 2564] = 1'b0;  addr_rom[ 2564]='h00000010;  wr_data_rom[ 2564]='h00000000;
    rd_cycle[ 2565] = 1'b1;  wr_cycle[ 2565] = 1'b0;  addr_rom[ 2565]='h00000014;  wr_data_rom[ 2565]='h00000000;
    rd_cycle[ 2566] = 1'b1;  wr_cycle[ 2566] = 1'b0;  addr_rom[ 2566]='h00000018;  wr_data_rom[ 2566]='h00000000;
    rd_cycle[ 2567] = 1'b1;  wr_cycle[ 2567] = 1'b0;  addr_rom[ 2567]='h0000001c;  wr_data_rom[ 2567]='h00000000;
    rd_cycle[ 2568] = 1'b1;  wr_cycle[ 2568] = 1'b0;  addr_rom[ 2568]='h00000020;  wr_data_rom[ 2568]='h00000000;
    rd_cycle[ 2569] = 1'b1;  wr_cycle[ 2569] = 1'b0;  addr_rom[ 2569]='h00000024;  wr_data_rom[ 2569]='h00000000;
    rd_cycle[ 2570] = 1'b1;  wr_cycle[ 2570] = 1'b0;  addr_rom[ 2570]='h00000028;  wr_data_rom[ 2570]='h00000000;
    rd_cycle[ 2571] = 1'b1;  wr_cycle[ 2571] = 1'b0;  addr_rom[ 2571]='h0000002c;  wr_data_rom[ 2571]='h00000000;
    rd_cycle[ 2572] = 1'b1;  wr_cycle[ 2572] = 1'b0;  addr_rom[ 2572]='h00000030;  wr_data_rom[ 2572]='h00000000;
    rd_cycle[ 2573] = 1'b1;  wr_cycle[ 2573] = 1'b0;  addr_rom[ 2573]='h00000034;  wr_data_rom[ 2573]='h00000000;
    rd_cycle[ 2574] = 1'b1;  wr_cycle[ 2574] = 1'b0;  addr_rom[ 2574]='h00000038;  wr_data_rom[ 2574]='h00000000;
    rd_cycle[ 2575] = 1'b1;  wr_cycle[ 2575] = 1'b0;  addr_rom[ 2575]='h0000003c;  wr_data_rom[ 2575]='h00000000;
    rd_cycle[ 2576] = 1'b1;  wr_cycle[ 2576] = 1'b0;  addr_rom[ 2576]='h00000040;  wr_data_rom[ 2576]='h00000000;
    rd_cycle[ 2577] = 1'b1;  wr_cycle[ 2577] = 1'b0;  addr_rom[ 2577]='h00000044;  wr_data_rom[ 2577]='h00000000;
    rd_cycle[ 2578] = 1'b1;  wr_cycle[ 2578] = 1'b0;  addr_rom[ 2578]='h00000048;  wr_data_rom[ 2578]='h00000000;
    rd_cycle[ 2579] = 1'b1;  wr_cycle[ 2579] = 1'b0;  addr_rom[ 2579]='h0000004c;  wr_data_rom[ 2579]='h00000000;
    rd_cycle[ 2580] = 1'b1;  wr_cycle[ 2580] = 1'b0;  addr_rom[ 2580]='h00000050;  wr_data_rom[ 2580]='h00000000;
    rd_cycle[ 2581] = 1'b1;  wr_cycle[ 2581] = 1'b0;  addr_rom[ 2581]='h00000054;  wr_data_rom[ 2581]='h00000000;
    rd_cycle[ 2582] = 1'b1;  wr_cycle[ 2582] = 1'b0;  addr_rom[ 2582]='h00000058;  wr_data_rom[ 2582]='h00000000;
    rd_cycle[ 2583] = 1'b1;  wr_cycle[ 2583] = 1'b0;  addr_rom[ 2583]='h0000005c;  wr_data_rom[ 2583]='h00000000;
    rd_cycle[ 2584] = 1'b1;  wr_cycle[ 2584] = 1'b0;  addr_rom[ 2584]='h00000060;  wr_data_rom[ 2584]='h00000000;
    rd_cycle[ 2585] = 1'b1;  wr_cycle[ 2585] = 1'b0;  addr_rom[ 2585]='h00000064;  wr_data_rom[ 2585]='h00000000;
    rd_cycle[ 2586] = 1'b1;  wr_cycle[ 2586] = 1'b0;  addr_rom[ 2586]='h00000068;  wr_data_rom[ 2586]='h00000000;
    rd_cycle[ 2587] = 1'b1;  wr_cycle[ 2587] = 1'b0;  addr_rom[ 2587]='h0000006c;  wr_data_rom[ 2587]='h00000000;
    rd_cycle[ 2588] = 1'b1;  wr_cycle[ 2588] = 1'b0;  addr_rom[ 2588]='h00000070;  wr_data_rom[ 2588]='h00000000;
    rd_cycle[ 2589] = 1'b1;  wr_cycle[ 2589] = 1'b0;  addr_rom[ 2589]='h00000074;  wr_data_rom[ 2589]='h00000000;
    rd_cycle[ 2590] = 1'b1;  wr_cycle[ 2590] = 1'b0;  addr_rom[ 2590]='h00000078;  wr_data_rom[ 2590]='h00000000;
    rd_cycle[ 2591] = 1'b1;  wr_cycle[ 2591] = 1'b0;  addr_rom[ 2591]='h0000007c;  wr_data_rom[ 2591]='h00000000;
    rd_cycle[ 2592] = 1'b1;  wr_cycle[ 2592] = 1'b0;  addr_rom[ 2592]='h00000080;  wr_data_rom[ 2592]='h00000000;
    rd_cycle[ 2593] = 1'b1;  wr_cycle[ 2593] = 1'b0;  addr_rom[ 2593]='h00000084;  wr_data_rom[ 2593]='h00000000;
    rd_cycle[ 2594] = 1'b1;  wr_cycle[ 2594] = 1'b0;  addr_rom[ 2594]='h00000088;  wr_data_rom[ 2594]='h00000000;
    rd_cycle[ 2595] = 1'b1;  wr_cycle[ 2595] = 1'b0;  addr_rom[ 2595]='h0000008c;  wr_data_rom[ 2595]='h00000000;
    rd_cycle[ 2596] = 1'b1;  wr_cycle[ 2596] = 1'b0;  addr_rom[ 2596]='h00000090;  wr_data_rom[ 2596]='h00000000;
    rd_cycle[ 2597] = 1'b1;  wr_cycle[ 2597] = 1'b0;  addr_rom[ 2597]='h00000094;  wr_data_rom[ 2597]='h00000000;
    rd_cycle[ 2598] = 1'b1;  wr_cycle[ 2598] = 1'b0;  addr_rom[ 2598]='h00000098;  wr_data_rom[ 2598]='h00000000;
    rd_cycle[ 2599] = 1'b1;  wr_cycle[ 2599] = 1'b0;  addr_rom[ 2599]='h0000009c;  wr_data_rom[ 2599]='h00000000;
    rd_cycle[ 2600] = 1'b1;  wr_cycle[ 2600] = 1'b0;  addr_rom[ 2600]='h000000a0;  wr_data_rom[ 2600]='h00000000;
    rd_cycle[ 2601] = 1'b1;  wr_cycle[ 2601] = 1'b0;  addr_rom[ 2601]='h000000a4;  wr_data_rom[ 2601]='h00000000;
    rd_cycle[ 2602] = 1'b1;  wr_cycle[ 2602] = 1'b0;  addr_rom[ 2602]='h000000a8;  wr_data_rom[ 2602]='h00000000;
    rd_cycle[ 2603] = 1'b1;  wr_cycle[ 2603] = 1'b0;  addr_rom[ 2603]='h000000ac;  wr_data_rom[ 2603]='h00000000;
    rd_cycle[ 2604] = 1'b1;  wr_cycle[ 2604] = 1'b0;  addr_rom[ 2604]='h000000b0;  wr_data_rom[ 2604]='h00000000;
    rd_cycle[ 2605] = 1'b1;  wr_cycle[ 2605] = 1'b0;  addr_rom[ 2605]='h000000b4;  wr_data_rom[ 2605]='h00000000;
    rd_cycle[ 2606] = 1'b1;  wr_cycle[ 2606] = 1'b0;  addr_rom[ 2606]='h000000b8;  wr_data_rom[ 2606]='h00000000;
    rd_cycle[ 2607] = 1'b1;  wr_cycle[ 2607] = 1'b0;  addr_rom[ 2607]='h000000bc;  wr_data_rom[ 2607]='h00000000;
    rd_cycle[ 2608] = 1'b1;  wr_cycle[ 2608] = 1'b0;  addr_rom[ 2608]='h000000c0;  wr_data_rom[ 2608]='h00000000;
    rd_cycle[ 2609] = 1'b1;  wr_cycle[ 2609] = 1'b0;  addr_rom[ 2609]='h000000c4;  wr_data_rom[ 2609]='h00000000;
    rd_cycle[ 2610] = 1'b1;  wr_cycle[ 2610] = 1'b0;  addr_rom[ 2610]='h000000c8;  wr_data_rom[ 2610]='h00000000;
    rd_cycle[ 2611] = 1'b1;  wr_cycle[ 2611] = 1'b0;  addr_rom[ 2611]='h000000cc;  wr_data_rom[ 2611]='h00000000;
    rd_cycle[ 2612] = 1'b1;  wr_cycle[ 2612] = 1'b0;  addr_rom[ 2612]='h000000d0;  wr_data_rom[ 2612]='h00000000;
    rd_cycle[ 2613] = 1'b1;  wr_cycle[ 2613] = 1'b0;  addr_rom[ 2613]='h000000d4;  wr_data_rom[ 2613]='h00000000;
    rd_cycle[ 2614] = 1'b1;  wr_cycle[ 2614] = 1'b0;  addr_rom[ 2614]='h000000d8;  wr_data_rom[ 2614]='h00000000;
    rd_cycle[ 2615] = 1'b1;  wr_cycle[ 2615] = 1'b0;  addr_rom[ 2615]='h000000dc;  wr_data_rom[ 2615]='h00000000;
    rd_cycle[ 2616] = 1'b1;  wr_cycle[ 2616] = 1'b0;  addr_rom[ 2616]='h000000e0;  wr_data_rom[ 2616]='h00000000;
    rd_cycle[ 2617] = 1'b1;  wr_cycle[ 2617] = 1'b0;  addr_rom[ 2617]='h000000e4;  wr_data_rom[ 2617]='h00000000;
    rd_cycle[ 2618] = 1'b1;  wr_cycle[ 2618] = 1'b0;  addr_rom[ 2618]='h000000e8;  wr_data_rom[ 2618]='h00000000;
    rd_cycle[ 2619] = 1'b1;  wr_cycle[ 2619] = 1'b0;  addr_rom[ 2619]='h000000ec;  wr_data_rom[ 2619]='h00000000;
    rd_cycle[ 2620] = 1'b1;  wr_cycle[ 2620] = 1'b0;  addr_rom[ 2620]='h000000f0;  wr_data_rom[ 2620]='h00000000;
    rd_cycle[ 2621] = 1'b1;  wr_cycle[ 2621] = 1'b0;  addr_rom[ 2621]='h000000f4;  wr_data_rom[ 2621]='h00000000;
    rd_cycle[ 2622] = 1'b1;  wr_cycle[ 2622] = 1'b0;  addr_rom[ 2622]='h000000f8;  wr_data_rom[ 2622]='h00000000;
    rd_cycle[ 2623] = 1'b1;  wr_cycle[ 2623] = 1'b0;  addr_rom[ 2623]='h000000fc;  wr_data_rom[ 2623]='h00000000;
    rd_cycle[ 2624] = 1'b1;  wr_cycle[ 2624] = 1'b0;  addr_rom[ 2624]='h00000100;  wr_data_rom[ 2624]='h00000000;
    rd_cycle[ 2625] = 1'b1;  wr_cycle[ 2625] = 1'b0;  addr_rom[ 2625]='h00000104;  wr_data_rom[ 2625]='h00000000;
    rd_cycle[ 2626] = 1'b1;  wr_cycle[ 2626] = 1'b0;  addr_rom[ 2626]='h00000108;  wr_data_rom[ 2626]='h00000000;
    rd_cycle[ 2627] = 1'b1;  wr_cycle[ 2627] = 1'b0;  addr_rom[ 2627]='h0000010c;  wr_data_rom[ 2627]='h00000000;
    rd_cycle[ 2628] = 1'b1;  wr_cycle[ 2628] = 1'b0;  addr_rom[ 2628]='h00000110;  wr_data_rom[ 2628]='h00000000;
    rd_cycle[ 2629] = 1'b1;  wr_cycle[ 2629] = 1'b0;  addr_rom[ 2629]='h00000114;  wr_data_rom[ 2629]='h00000000;
    rd_cycle[ 2630] = 1'b1;  wr_cycle[ 2630] = 1'b0;  addr_rom[ 2630]='h00000118;  wr_data_rom[ 2630]='h00000000;
    rd_cycle[ 2631] = 1'b1;  wr_cycle[ 2631] = 1'b0;  addr_rom[ 2631]='h0000011c;  wr_data_rom[ 2631]='h00000000;
    rd_cycle[ 2632] = 1'b1;  wr_cycle[ 2632] = 1'b0;  addr_rom[ 2632]='h00000120;  wr_data_rom[ 2632]='h00000000;
    rd_cycle[ 2633] = 1'b1;  wr_cycle[ 2633] = 1'b0;  addr_rom[ 2633]='h00000124;  wr_data_rom[ 2633]='h00000000;
    rd_cycle[ 2634] = 1'b1;  wr_cycle[ 2634] = 1'b0;  addr_rom[ 2634]='h00000128;  wr_data_rom[ 2634]='h00000000;
    rd_cycle[ 2635] = 1'b1;  wr_cycle[ 2635] = 1'b0;  addr_rom[ 2635]='h0000012c;  wr_data_rom[ 2635]='h00000000;
    rd_cycle[ 2636] = 1'b1;  wr_cycle[ 2636] = 1'b0;  addr_rom[ 2636]='h00000130;  wr_data_rom[ 2636]='h00000000;
    rd_cycle[ 2637] = 1'b1;  wr_cycle[ 2637] = 1'b0;  addr_rom[ 2637]='h00000134;  wr_data_rom[ 2637]='h00000000;
    rd_cycle[ 2638] = 1'b1;  wr_cycle[ 2638] = 1'b0;  addr_rom[ 2638]='h00000138;  wr_data_rom[ 2638]='h00000000;
    rd_cycle[ 2639] = 1'b1;  wr_cycle[ 2639] = 1'b0;  addr_rom[ 2639]='h0000013c;  wr_data_rom[ 2639]='h00000000;
    rd_cycle[ 2640] = 1'b1;  wr_cycle[ 2640] = 1'b0;  addr_rom[ 2640]='h00000140;  wr_data_rom[ 2640]='h00000000;
    rd_cycle[ 2641] = 1'b1;  wr_cycle[ 2641] = 1'b0;  addr_rom[ 2641]='h00000144;  wr_data_rom[ 2641]='h00000000;
    rd_cycle[ 2642] = 1'b1;  wr_cycle[ 2642] = 1'b0;  addr_rom[ 2642]='h00000148;  wr_data_rom[ 2642]='h00000000;
    rd_cycle[ 2643] = 1'b1;  wr_cycle[ 2643] = 1'b0;  addr_rom[ 2643]='h0000014c;  wr_data_rom[ 2643]='h00000000;
    rd_cycle[ 2644] = 1'b1;  wr_cycle[ 2644] = 1'b0;  addr_rom[ 2644]='h00000150;  wr_data_rom[ 2644]='h00000000;
    rd_cycle[ 2645] = 1'b1;  wr_cycle[ 2645] = 1'b0;  addr_rom[ 2645]='h00000154;  wr_data_rom[ 2645]='h00000000;
    rd_cycle[ 2646] = 1'b1;  wr_cycle[ 2646] = 1'b0;  addr_rom[ 2646]='h00000158;  wr_data_rom[ 2646]='h00000000;
    rd_cycle[ 2647] = 1'b1;  wr_cycle[ 2647] = 1'b0;  addr_rom[ 2647]='h0000015c;  wr_data_rom[ 2647]='h00000000;
    rd_cycle[ 2648] = 1'b1;  wr_cycle[ 2648] = 1'b0;  addr_rom[ 2648]='h00000160;  wr_data_rom[ 2648]='h00000000;
    rd_cycle[ 2649] = 1'b1;  wr_cycle[ 2649] = 1'b0;  addr_rom[ 2649]='h00000164;  wr_data_rom[ 2649]='h00000000;
    rd_cycle[ 2650] = 1'b1;  wr_cycle[ 2650] = 1'b0;  addr_rom[ 2650]='h00000168;  wr_data_rom[ 2650]='h00000000;
    rd_cycle[ 2651] = 1'b1;  wr_cycle[ 2651] = 1'b0;  addr_rom[ 2651]='h0000016c;  wr_data_rom[ 2651]='h00000000;
    rd_cycle[ 2652] = 1'b1;  wr_cycle[ 2652] = 1'b0;  addr_rom[ 2652]='h00000170;  wr_data_rom[ 2652]='h00000000;
    rd_cycle[ 2653] = 1'b1;  wr_cycle[ 2653] = 1'b0;  addr_rom[ 2653]='h00000174;  wr_data_rom[ 2653]='h00000000;
    rd_cycle[ 2654] = 1'b1;  wr_cycle[ 2654] = 1'b0;  addr_rom[ 2654]='h00000178;  wr_data_rom[ 2654]='h00000000;
    rd_cycle[ 2655] = 1'b1;  wr_cycle[ 2655] = 1'b0;  addr_rom[ 2655]='h0000017c;  wr_data_rom[ 2655]='h00000000;
    rd_cycle[ 2656] = 1'b1;  wr_cycle[ 2656] = 1'b0;  addr_rom[ 2656]='h00000180;  wr_data_rom[ 2656]='h00000000;
    rd_cycle[ 2657] = 1'b1;  wr_cycle[ 2657] = 1'b0;  addr_rom[ 2657]='h00000184;  wr_data_rom[ 2657]='h00000000;
    rd_cycle[ 2658] = 1'b1;  wr_cycle[ 2658] = 1'b0;  addr_rom[ 2658]='h00000188;  wr_data_rom[ 2658]='h00000000;
    rd_cycle[ 2659] = 1'b1;  wr_cycle[ 2659] = 1'b0;  addr_rom[ 2659]='h0000018c;  wr_data_rom[ 2659]='h00000000;
    rd_cycle[ 2660] = 1'b1;  wr_cycle[ 2660] = 1'b0;  addr_rom[ 2660]='h00000190;  wr_data_rom[ 2660]='h00000000;
    rd_cycle[ 2661] = 1'b1;  wr_cycle[ 2661] = 1'b0;  addr_rom[ 2661]='h00000194;  wr_data_rom[ 2661]='h00000000;
    rd_cycle[ 2662] = 1'b1;  wr_cycle[ 2662] = 1'b0;  addr_rom[ 2662]='h00000198;  wr_data_rom[ 2662]='h00000000;
    rd_cycle[ 2663] = 1'b1;  wr_cycle[ 2663] = 1'b0;  addr_rom[ 2663]='h0000019c;  wr_data_rom[ 2663]='h00000000;
    rd_cycle[ 2664] = 1'b1;  wr_cycle[ 2664] = 1'b0;  addr_rom[ 2664]='h000001a0;  wr_data_rom[ 2664]='h00000000;
    rd_cycle[ 2665] = 1'b1;  wr_cycle[ 2665] = 1'b0;  addr_rom[ 2665]='h000001a4;  wr_data_rom[ 2665]='h00000000;
    rd_cycle[ 2666] = 1'b1;  wr_cycle[ 2666] = 1'b0;  addr_rom[ 2666]='h000001a8;  wr_data_rom[ 2666]='h00000000;
    rd_cycle[ 2667] = 1'b1;  wr_cycle[ 2667] = 1'b0;  addr_rom[ 2667]='h000001ac;  wr_data_rom[ 2667]='h00000000;
    rd_cycle[ 2668] = 1'b1;  wr_cycle[ 2668] = 1'b0;  addr_rom[ 2668]='h000001b0;  wr_data_rom[ 2668]='h00000000;
    rd_cycle[ 2669] = 1'b1;  wr_cycle[ 2669] = 1'b0;  addr_rom[ 2669]='h000001b4;  wr_data_rom[ 2669]='h00000000;
    rd_cycle[ 2670] = 1'b1;  wr_cycle[ 2670] = 1'b0;  addr_rom[ 2670]='h000001b8;  wr_data_rom[ 2670]='h00000000;
    rd_cycle[ 2671] = 1'b1;  wr_cycle[ 2671] = 1'b0;  addr_rom[ 2671]='h000001bc;  wr_data_rom[ 2671]='h00000000;
    rd_cycle[ 2672] = 1'b1;  wr_cycle[ 2672] = 1'b0;  addr_rom[ 2672]='h000001c0;  wr_data_rom[ 2672]='h00000000;
    rd_cycle[ 2673] = 1'b1;  wr_cycle[ 2673] = 1'b0;  addr_rom[ 2673]='h000001c4;  wr_data_rom[ 2673]='h00000000;
    rd_cycle[ 2674] = 1'b1;  wr_cycle[ 2674] = 1'b0;  addr_rom[ 2674]='h000001c8;  wr_data_rom[ 2674]='h00000000;
    rd_cycle[ 2675] = 1'b1;  wr_cycle[ 2675] = 1'b0;  addr_rom[ 2675]='h000001cc;  wr_data_rom[ 2675]='h00000000;
    rd_cycle[ 2676] = 1'b1;  wr_cycle[ 2676] = 1'b0;  addr_rom[ 2676]='h000001d0;  wr_data_rom[ 2676]='h00000000;
    rd_cycle[ 2677] = 1'b1;  wr_cycle[ 2677] = 1'b0;  addr_rom[ 2677]='h000001d4;  wr_data_rom[ 2677]='h00000000;
    rd_cycle[ 2678] = 1'b1;  wr_cycle[ 2678] = 1'b0;  addr_rom[ 2678]='h000001d8;  wr_data_rom[ 2678]='h00000000;
    rd_cycle[ 2679] = 1'b1;  wr_cycle[ 2679] = 1'b0;  addr_rom[ 2679]='h000001dc;  wr_data_rom[ 2679]='h00000000;
    rd_cycle[ 2680] = 1'b1;  wr_cycle[ 2680] = 1'b0;  addr_rom[ 2680]='h000001e0;  wr_data_rom[ 2680]='h00000000;
    rd_cycle[ 2681] = 1'b1;  wr_cycle[ 2681] = 1'b0;  addr_rom[ 2681]='h000001e4;  wr_data_rom[ 2681]='h00000000;
    rd_cycle[ 2682] = 1'b1;  wr_cycle[ 2682] = 1'b0;  addr_rom[ 2682]='h000001e8;  wr_data_rom[ 2682]='h00000000;
    rd_cycle[ 2683] = 1'b1;  wr_cycle[ 2683] = 1'b0;  addr_rom[ 2683]='h000001ec;  wr_data_rom[ 2683]='h00000000;
    rd_cycle[ 2684] = 1'b1;  wr_cycle[ 2684] = 1'b0;  addr_rom[ 2684]='h000001f0;  wr_data_rom[ 2684]='h00000000;
    rd_cycle[ 2685] = 1'b1;  wr_cycle[ 2685] = 1'b0;  addr_rom[ 2685]='h000001f4;  wr_data_rom[ 2685]='h00000000;
    rd_cycle[ 2686] = 1'b1;  wr_cycle[ 2686] = 1'b0;  addr_rom[ 2686]='h000001f8;  wr_data_rom[ 2686]='h00000000;
    rd_cycle[ 2687] = 1'b1;  wr_cycle[ 2687] = 1'b0;  addr_rom[ 2687]='h000001fc;  wr_data_rom[ 2687]='h00000000;
    rd_cycle[ 2688] = 1'b1;  wr_cycle[ 2688] = 1'b0;  addr_rom[ 2688]='h00000200;  wr_data_rom[ 2688]='h00000000;
    rd_cycle[ 2689] = 1'b1;  wr_cycle[ 2689] = 1'b0;  addr_rom[ 2689]='h00000204;  wr_data_rom[ 2689]='h00000000;
    rd_cycle[ 2690] = 1'b1;  wr_cycle[ 2690] = 1'b0;  addr_rom[ 2690]='h00000208;  wr_data_rom[ 2690]='h00000000;
    rd_cycle[ 2691] = 1'b1;  wr_cycle[ 2691] = 1'b0;  addr_rom[ 2691]='h0000020c;  wr_data_rom[ 2691]='h00000000;
    rd_cycle[ 2692] = 1'b1;  wr_cycle[ 2692] = 1'b0;  addr_rom[ 2692]='h00000210;  wr_data_rom[ 2692]='h00000000;
    rd_cycle[ 2693] = 1'b1;  wr_cycle[ 2693] = 1'b0;  addr_rom[ 2693]='h00000214;  wr_data_rom[ 2693]='h00000000;
    rd_cycle[ 2694] = 1'b1;  wr_cycle[ 2694] = 1'b0;  addr_rom[ 2694]='h00000218;  wr_data_rom[ 2694]='h00000000;
    rd_cycle[ 2695] = 1'b1;  wr_cycle[ 2695] = 1'b0;  addr_rom[ 2695]='h0000021c;  wr_data_rom[ 2695]='h00000000;
    rd_cycle[ 2696] = 1'b1;  wr_cycle[ 2696] = 1'b0;  addr_rom[ 2696]='h00000220;  wr_data_rom[ 2696]='h00000000;
    rd_cycle[ 2697] = 1'b1;  wr_cycle[ 2697] = 1'b0;  addr_rom[ 2697]='h00000224;  wr_data_rom[ 2697]='h00000000;
    rd_cycle[ 2698] = 1'b1;  wr_cycle[ 2698] = 1'b0;  addr_rom[ 2698]='h00000228;  wr_data_rom[ 2698]='h00000000;
    rd_cycle[ 2699] = 1'b1;  wr_cycle[ 2699] = 1'b0;  addr_rom[ 2699]='h0000022c;  wr_data_rom[ 2699]='h00000000;
    rd_cycle[ 2700] = 1'b1;  wr_cycle[ 2700] = 1'b0;  addr_rom[ 2700]='h00000230;  wr_data_rom[ 2700]='h00000000;
    rd_cycle[ 2701] = 1'b1;  wr_cycle[ 2701] = 1'b0;  addr_rom[ 2701]='h00000234;  wr_data_rom[ 2701]='h00000000;
    rd_cycle[ 2702] = 1'b1;  wr_cycle[ 2702] = 1'b0;  addr_rom[ 2702]='h00000238;  wr_data_rom[ 2702]='h00000000;
    rd_cycle[ 2703] = 1'b1;  wr_cycle[ 2703] = 1'b0;  addr_rom[ 2703]='h0000023c;  wr_data_rom[ 2703]='h00000000;
    rd_cycle[ 2704] = 1'b1;  wr_cycle[ 2704] = 1'b0;  addr_rom[ 2704]='h00000240;  wr_data_rom[ 2704]='h00000000;
    rd_cycle[ 2705] = 1'b1;  wr_cycle[ 2705] = 1'b0;  addr_rom[ 2705]='h00000244;  wr_data_rom[ 2705]='h00000000;
    rd_cycle[ 2706] = 1'b1;  wr_cycle[ 2706] = 1'b0;  addr_rom[ 2706]='h00000248;  wr_data_rom[ 2706]='h00000000;
    rd_cycle[ 2707] = 1'b1;  wr_cycle[ 2707] = 1'b0;  addr_rom[ 2707]='h0000024c;  wr_data_rom[ 2707]='h00000000;
    rd_cycle[ 2708] = 1'b1;  wr_cycle[ 2708] = 1'b0;  addr_rom[ 2708]='h00000250;  wr_data_rom[ 2708]='h00000000;
    rd_cycle[ 2709] = 1'b1;  wr_cycle[ 2709] = 1'b0;  addr_rom[ 2709]='h00000254;  wr_data_rom[ 2709]='h00000000;
    rd_cycle[ 2710] = 1'b1;  wr_cycle[ 2710] = 1'b0;  addr_rom[ 2710]='h00000258;  wr_data_rom[ 2710]='h00000000;
    rd_cycle[ 2711] = 1'b1;  wr_cycle[ 2711] = 1'b0;  addr_rom[ 2711]='h0000025c;  wr_data_rom[ 2711]='h00000000;
    rd_cycle[ 2712] = 1'b1;  wr_cycle[ 2712] = 1'b0;  addr_rom[ 2712]='h00000260;  wr_data_rom[ 2712]='h00000000;
    rd_cycle[ 2713] = 1'b1;  wr_cycle[ 2713] = 1'b0;  addr_rom[ 2713]='h00000264;  wr_data_rom[ 2713]='h00000000;
    rd_cycle[ 2714] = 1'b1;  wr_cycle[ 2714] = 1'b0;  addr_rom[ 2714]='h00000268;  wr_data_rom[ 2714]='h00000000;
    rd_cycle[ 2715] = 1'b1;  wr_cycle[ 2715] = 1'b0;  addr_rom[ 2715]='h0000026c;  wr_data_rom[ 2715]='h00000000;
    rd_cycle[ 2716] = 1'b1;  wr_cycle[ 2716] = 1'b0;  addr_rom[ 2716]='h00000270;  wr_data_rom[ 2716]='h00000000;
    rd_cycle[ 2717] = 1'b1;  wr_cycle[ 2717] = 1'b0;  addr_rom[ 2717]='h00000274;  wr_data_rom[ 2717]='h00000000;
    rd_cycle[ 2718] = 1'b1;  wr_cycle[ 2718] = 1'b0;  addr_rom[ 2718]='h00000278;  wr_data_rom[ 2718]='h00000000;
    rd_cycle[ 2719] = 1'b1;  wr_cycle[ 2719] = 1'b0;  addr_rom[ 2719]='h0000027c;  wr_data_rom[ 2719]='h00000000;
    rd_cycle[ 2720] = 1'b1;  wr_cycle[ 2720] = 1'b0;  addr_rom[ 2720]='h00000280;  wr_data_rom[ 2720]='h00000000;
    rd_cycle[ 2721] = 1'b1;  wr_cycle[ 2721] = 1'b0;  addr_rom[ 2721]='h00000284;  wr_data_rom[ 2721]='h00000000;
    rd_cycle[ 2722] = 1'b1;  wr_cycle[ 2722] = 1'b0;  addr_rom[ 2722]='h00000288;  wr_data_rom[ 2722]='h00000000;
    rd_cycle[ 2723] = 1'b1;  wr_cycle[ 2723] = 1'b0;  addr_rom[ 2723]='h0000028c;  wr_data_rom[ 2723]='h00000000;
    rd_cycle[ 2724] = 1'b1;  wr_cycle[ 2724] = 1'b0;  addr_rom[ 2724]='h00000290;  wr_data_rom[ 2724]='h00000000;
    rd_cycle[ 2725] = 1'b1;  wr_cycle[ 2725] = 1'b0;  addr_rom[ 2725]='h00000294;  wr_data_rom[ 2725]='h00000000;
    rd_cycle[ 2726] = 1'b1;  wr_cycle[ 2726] = 1'b0;  addr_rom[ 2726]='h00000298;  wr_data_rom[ 2726]='h00000000;
    rd_cycle[ 2727] = 1'b1;  wr_cycle[ 2727] = 1'b0;  addr_rom[ 2727]='h0000029c;  wr_data_rom[ 2727]='h00000000;
    rd_cycle[ 2728] = 1'b1;  wr_cycle[ 2728] = 1'b0;  addr_rom[ 2728]='h000002a0;  wr_data_rom[ 2728]='h00000000;
    rd_cycle[ 2729] = 1'b1;  wr_cycle[ 2729] = 1'b0;  addr_rom[ 2729]='h000002a4;  wr_data_rom[ 2729]='h00000000;
    rd_cycle[ 2730] = 1'b1;  wr_cycle[ 2730] = 1'b0;  addr_rom[ 2730]='h000002a8;  wr_data_rom[ 2730]='h00000000;
    rd_cycle[ 2731] = 1'b1;  wr_cycle[ 2731] = 1'b0;  addr_rom[ 2731]='h000002ac;  wr_data_rom[ 2731]='h00000000;
    rd_cycle[ 2732] = 1'b1;  wr_cycle[ 2732] = 1'b0;  addr_rom[ 2732]='h000002b0;  wr_data_rom[ 2732]='h00000000;
    rd_cycle[ 2733] = 1'b1;  wr_cycle[ 2733] = 1'b0;  addr_rom[ 2733]='h000002b4;  wr_data_rom[ 2733]='h00000000;
    rd_cycle[ 2734] = 1'b1;  wr_cycle[ 2734] = 1'b0;  addr_rom[ 2734]='h000002b8;  wr_data_rom[ 2734]='h00000000;
    rd_cycle[ 2735] = 1'b1;  wr_cycle[ 2735] = 1'b0;  addr_rom[ 2735]='h000002bc;  wr_data_rom[ 2735]='h00000000;
    rd_cycle[ 2736] = 1'b1;  wr_cycle[ 2736] = 1'b0;  addr_rom[ 2736]='h000002c0;  wr_data_rom[ 2736]='h00000000;
    rd_cycle[ 2737] = 1'b1;  wr_cycle[ 2737] = 1'b0;  addr_rom[ 2737]='h000002c4;  wr_data_rom[ 2737]='h00000000;
    rd_cycle[ 2738] = 1'b1;  wr_cycle[ 2738] = 1'b0;  addr_rom[ 2738]='h000002c8;  wr_data_rom[ 2738]='h00000000;
    rd_cycle[ 2739] = 1'b1;  wr_cycle[ 2739] = 1'b0;  addr_rom[ 2739]='h000002cc;  wr_data_rom[ 2739]='h00000000;
    rd_cycle[ 2740] = 1'b1;  wr_cycle[ 2740] = 1'b0;  addr_rom[ 2740]='h000002d0;  wr_data_rom[ 2740]='h00000000;
    rd_cycle[ 2741] = 1'b1;  wr_cycle[ 2741] = 1'b0;  addr_rom[ 2741]='h000002d4;  wr_data_rom[ 2741]='h00000000;
    rd_cycle[ 2742] = 1'b1;  wr_cycle[ 2742] = 1'b0;  addr_rom[ 2742]='h000002d8;  wr_data_rom[ 2742]='h00000000;
    rd_cycle[ 2743] = 1'b1;  wr_cycle[ 2743] = 1'b0;  addr_rom[ 2743]='h000002dc;  wr_data_rom[ 2743]='h00000000;
    rd_cycle[ 2744] = 1'b1;  wr_cycle[ 2744] = 1'b0;  addr_rom[ 2744]='h000002e0;  wr_data_rom[ 2744]='h00000000;
    rd_cycle[ 2745] = 1'b1;  wr_cycle[ 2745] = 1'b0;  addr_rom[ 2745]='h000002e4;  wr_data_rom[ 2745]='h00000000;
    rd_cycle[ 2746] = 1'b1;  wr_cycle[ 2746] = 1'b0;  addr_rom[ 2746]='h000002e8;  wr_data_rom[ 2746]='h00000000;
    rd_cycle[ 2747] = 1'b1;  wr_cycle[ 2747] = 1'b0;  addr_rom[ 2747]='h000002ec;  wr_data_rom[ 2747]='h00000000;
    rd_cycle[ 2748] = 1'b1;  wr_cycle[ 2748] = 1'b0;  addr_rom[ 2748]='h000002f0;  wr_data_rom[ 2748]='h00000000;
    rd_cycle[ 2749] = 1'b1;  wr_cycle[ 2749] = 1'b0;  addr_rom[ 2749]='h000002f4;  wr_data_rom[ 2749]='h00000000;
    rd_cycle[ 2750] = 1'b1;  wr_cycle[ 2750] = 1'b0;  addr_rom[ 2750]='h000002f8;  wr_data_rom[ 2750]='h00000000;
    rd_cycle[ 2751] = 1'b1;  wr_cycle[ 2751] = 1'b0;  addr_rom[ 2751]='h000002fc;  wr_data_rom[ 2751]='h00000000;
    rd_cycle[ 2752] = 1'b1;  wr_cycle[ 2752] = 1'b0;  addr_rom[ 2752]='h00000300;  wr_data_rom[ 2752]='h00000000;
    rd_cycle[ 2753] = 1'b1;  wr_cycle[ 2753] = 1'b0;  addr_rom[ 2753]='h00000304;  wr_data_rom[ 2753]='h00000000;
    rd_cycle[ 2754] = 1'b1;  wr_cycle[ 2754] = 1'b0;  addr_rom[ 2754]='h00000308;  wr_data_rom[ 2754]='h00000000;
    rd_cycle[ 2755] = 1'b1;  wr_cycle[ 2755] = 1'b0;  addr_rom[ 2755]='h0000030c;  wr_data_rom[ 2755]='h00000000;
    rd_cycle[ 2756] = 1'b1;  wr_cycle[ 2756] = 1'b0;  addr_rom[ 2756]='h00000310;  wr_data_rom[ 2756]='h00000000;
    rd_cycle[ 2757] = 1'b1;  wr_cycle[ 2757] = 1'b0;  addr_rom[ 2757]='h00000314;  wr_data_rom[ 2757]='h00000000;
    rd_cycle[ 2758] = 1'b1;  wr_cycle[ 2758] = 1'b0;  addr_rom[ 2758]='h00000318;  wr_data_rom[ 2758]='h00000000;
    rd_cycle[ 2759] = 1'b1;  wr_cycle[ 2759] = 1'b0;  addr_rom[ 2759]='h0000031c;  wr_data_rom[ 2759]='h00000000;
    rd_cycle[ 2760] = 1'b1;  wr_cycle[ 2760] = 1'b0;  addr_rom[ 2760]='h00000320;  wr_data_rom[ 2760]='h00000000;
    rd_cycle[ 2761] = 1'b1;  wr_cycle[ 2761] = 1'b0;  addr_rom[ 2761]='h00000324;  wr_data_rom[ 2761]='h00000000;
    rd_cycle[ 2762] = 1'b1;  wr_cycle[ 2762] = 1'b0;  addr_rom[ 2762]='h00000328;  wr_data_rom[ 2762]='h00000000;
    rd_cycle[ 2763] = 1'b1;  wr_cycle[ 2763] = 1'b0;  addr_rom[ 2763]='h0000032c;  wr_data_rom[ 2763]='h00000000;
    rd_cycle[ 2764] = 1'b1;  wr_cycle[ 2764] = 1'b0;  addr_rom[ 2764]='h00000330;  wr_data_rom[ 2764]='h00000000;
    rd_cycle[ 2765] = 1'b1;  wr_cycle[ 2765] = 1'b0;  addr_rom[ 2765]='h00000334;  wr_data_rom[ 2765]='h00000000;
    rd_cycle[ 2766] = 1'b1;  wr_cycle[ 2766] = 1'b0;  addr_rom[ 2766]='h00000338;  wr_data_rom[ 2766]='h00000000;
    rd_cycle[ 2767] = 1'b1;  wr_cycle[ 2767] = 1'b0;  addr_rom[ 2767]='h0000033c;  wr_data_rom[ 2767]='h00000000;
    rd_cycle[ 2768] = 1'b1;  wr_cycle[ 2768] = 1'b0;  addr_rom[ 2768]='h00000340;  wr_data_rom[ 2768]='h00000000;
    rd_cycle[ 2769] = 1'b1;  wr_cycle[ 2769] = 1'b0;  addr_rom[ 2769]='h00000344;  wr_data_rom[ 2769]='h00000000;
    rd_cycle[ 2770] = 1'b1;  wr_cycle[ 2770] = 1'b0;  addr_rom[ 2770]='h00000348;  wr_data_rom[ 2770]='h00000000;
    rd_cycle[ 2771] = 1'b1;  wr_cycle[ 2771] = 1'b0;  addr_rom[ 2771]='h0000034c;  wr_data_rom[ 2771]='h00000000;
    rd_cycle[ 2772] = 1'b1;  wr_cycle[ 2772] = 1'b0;  addr_rom[ 2772]='h00000350;  wr_data_rom[ 2772]='h00000000;
    rd_cycle[ 2773] = 1'b1;  wr_cycle[ 2773] = 1'b0;  addr_rom[ 2773]='h00000354;  wr_data_rom[ 2773]='h00000000;
    rd_cycle[ 2774] = 1'b1;  wr_cycle[ 2774] = 1'b0;  addr_rom[ 2774]='h00000358;  wr_data_rom[ 2774]='h00000000;
    rd_cycle[ 2775] = 1'b1;  wr_cycle[ 2775] = 1'b0;  addr_rom[ 2775]='h0000035c;  wr_data_rom[ 2775]='h00000000;
    rd_cycle[ 2776] = 1'b1;  wr_cycle[ 2776] = 1'b0;  addr_rom[ 2776]='h00000360;  wr_data_rom[ 2776]='h00000000;
    rd_cycle[ 2777] = 1'b1;  wr_cycle[ 2777] = 1'b0;  addr_rom[ 2777]='h00000364;  wr_data_rom[ 2777]='h00000000;
    rd_cycle[ 2778] = 1'b1;  wr_cycle[ 2778] = 1'b0;  addr_rom[ 2778]='h00000368;  wr_data_rom[ 2778]='h00000000;
    rd_cycle[ 2779] = 1'b1;  wr_cycle[ 2779] = 1'b0;  addr_rom[ 2779]='h0000036c;  wr_data_rom[ 2779]='h00000000;
    rd_cycle[ 2780] = 1'b1;  wr_cycle[ 2780] = 1'b0;  addr_rom[ 2780]='h00000370;  wr_data_rom[ 2780]='h00000000;
    rd_cycle[ 2781] = 1'b1;  wr_cycle[ 2781] = 1'b0;  addr_rom[ 2781]='h00000374;  wr_data_rom[ 2781]='h00000000;
    rd_cycle[ 2782] = 1'b1;  wr_cycle[ 2782] = 1'b0;  addr_rom[ 2782]='h00000378;  wr_data_rom[ 2782]='h00000000;
    rd_cycle[ 2783] = 1'b1;  wr_cycle[ 2783] = 1'b0;  addr_rom[ 2783]='h0000037c;  wr_data_rom[ 2783]='h00000000;
    rd_cycle[ 2784] = 1'b1;  wr_cycle[ 2784] = 1'b0;  addr_rom[ 2784]='h00000380;  wr_data_rom[ 2784]='h00000000;
    rd_cycle[ 2785] = 1'b1;  wr_cycle[ 2785] = 1'b0;  addr_rom[ 2785]='h00000384;  wr_data_rom[ 2785]='h00000000;
    rd_cycle[ 2786] = 1'b1;  wr_cycle[ 2786] = 1'b0;  addr_rom[ 2786]='h00000388;  wr_data_rom[ 2786]='h00000000;
    rd_cycle[ 2787] = 1'b1;  wr_cycle[ 2787] = 1'b0;  addr_rom[ 2787]='h0000038c;  wr_data_rom[ 2787]='h00000000;
    rd_cycle[ 2788] = 1'b1;  wr_cycle[ 2788] = 1'b0;  addr_rom[ 2788]='h00000390;  wr_data_rom[ 2788]='h00000000;
    rd_cycle[ 2789] = 1'b1;  wr_cycle[ 2789] = 1'b0;  addr_rom[ 2789]='h00000394;  wr_data_rom[ 2789]='h00000000;
    rd_cycle[ 2790] = 1'b1;  wr_cycle[ 2790] = 1'b0;  addr_rom[ 2790]='h00000398;  wr_data_rom[ 2790]='h00000000;
    rd_cycle[ 2791] = 1'b1;  wr_cycle[ 2791] = 1'b0;  addr_rom[ 2791]='h0000039c;  wr_data_rom[ 2791]='h00000000;
    rd_cycle[ 2792] = 1'b1;  wr_cycle[ 2792] = 1'b0;  addr_rom[ 2792]='h000003a0;  wr_data_rom[ 2792]='h00000000;
    rd_cycle[ 2793] = 1'b1;  wr_cycle[ 2793] = 1'b0;  addr_rom[ 2793]='h000003a4;  wr_data_rom[ 2793]='h00000000;
    rd_cycle[ 2794] = 1'b1;  wr_cycle[ 2794] = 1'b0;  addr_rom[ 2794]='h000003a8;  wr_data_rom[ 2794]='h00000000;
    rd_cycle[ 2795] = 1'b1;  wr_cycle[ 2795] = 1'b0;  addr_rom[ 2795]='h000003ac;  wr_data_rom[ 2795]='h00000000;
    rd_cycle[ 2796] = 1'b1;  wr_cycle[ 2796] = 1'b0;  addr_rom[ 2796]='h000003b0;  wr_data_rom[ 2796]='h00000000;
    rd_cycle[ 2797] = 1'b1;  wr_cycle[ 2797] = 1'b0;  addr_rom[ 2797]='h000003b4;  wr_data_rom[ 2797]='h00000000;
    rd_cycle[ 2798] = 1'b1;  wr_cycle[ 2798] = 1'b0;  addr_rom[ 2798]='h000003b8;  wr_data_rom[ 2798]='h00000000;
    rd_cycle[ 2799] = 1'b1;  wr_cycle[ 2799] = 1'b0;  addr_rom[ 2799]='h000003bc;  wr_data_rom[ 2799]='h00000000;
    rd_cycle[ 2800] = 1'b1;  wr_cycle[ 2800] = 1'b0;  addr_rom[ 2800]='h000003c0;  wr_data_rom[ 2800]='h00000000;
    rd_cycle[ 2801] = 1'b1;  wr_cycle[ 2801] = 1'b0;  addr_rom[ 2801]='h000003c4;  wr_data_rom[ 2801]='h00000000;
    rd_cycle[ 2802] = 1'b1;  wr_cycle[ 2802] = 1'b0;  addr_rom[ 2802]='h000003c8;  wr_data_rom[ 2802]='h00000000;
    rd_cycle[ 2803] = 1'b1;  wr_cycle[ 2803] = 1'b0;  addr_rom[ 2803]='h000003cc;  wr_data_rom[ 2803]='h00000000;
    rd_cycle[ 2804] = 1'b1;  wr_cycle[ 2804] = 1'b0;  addr_rom[ 2804]='h000003d0;  wr_data_rom[ 2804]='h00000000;
    rd_cycle[ 2805] = 1'b1;  wr_cycle[ 2805] = 1'b0;  addr_rom[ 2805]='h000003d4;  wr_data_rom[ 2805]='h00000000;
    rd_cycle[ 2806] = 1'b1;  wr_cycle[ 2806] = 1'b0;  addr_rom[ 2806]='h000003d8;  wr_data_rom[ 2806]='h00000000;
    rd_cycle[ 2807] = 1'b1;  wr_cycle[ 2807] = 1'b0;  addr_rom[ 2807]='h000003dc;  wr_data_rom[ 2807]='h00000000;
    rd_cycle[ 2808] = 1'b1;  wr_cycle[ 2808] = 1'b0;  addr_rom[ 2808]='h000003e0;  wr_data_rom[ 2808]='h00000000;
    rd_cycle[ 2809] = 1'b1;  wr_cycle[ 2809] = 1'b0;  addr_rom[ 2809]='h000003e4;  wr_data_rom[ 2809]='h00000000;
    rd_cycle[ 2810] = 1'b1;  wr_cycle[ 2810] = 1'b0;  addr_rom[ 2810]='h000003e8;  wr_data_rom[ 2810]='h00000000;
    rd_cycle[ 2811] = 1'b1;  wr_cycle[ 2811] = 1'b0;  addr_rom[ 2811]='h000003ec;  wr_data_rom[ 2811]='h00000000;
    rd_cycle[ 2812] = 1'b1;  wr_cycle[ 2812] = 1'b0;  addr_rom[ 2812]='h000003f0;  wr_data_rom[ 2812]='h00000000;
    rd_cycle[ 2813] = 1'b1;  wr_cycle[ 2813] = 1'b0;  addr_rom[ 2813]='h000003f4;  wr_data_rom[ 2813]='h00000000;
    rd_cycle[ 2814] = 1'b1;  wr_cycle[ 2814] = 1'b0;  addr_rom[ 2814]='h000003f8;  wr_data_rom[ 2814]='h00000000;
    rd_cycle[ 2815] = 1'b1;  wr_cycle[ 2815] = 1'b0;  addr_rom[ 2815]='h000003fc;  wr_data_rom[ 2815]='h00000000;
    rd_cycle[ 2816] = 1'b1;  wr_cycle[ 2816] = 1'b0;  addr_rom[ 2816]='h00000400;  wr_data_rom[ 2816]='h00000000;
    rd_cycle[ 2817] = 1'b1;  wr_cycle[ 2817] = 1'b0;  addr_rom[ 2817]='h00000404;  wr_data_rom[ 2817]='h00000000;
    rd_cycle[ 2818] = 1'b1;  wr_cycle[ 2818] = 1'b0;  addr_rom[ 2818]='h00000408;  wr_data_rom[ 2818]='h00000000;
    rd_cycle[ 2819] = 1'b1;  wr_cycle[ 2819] = 1'b0;  addr_rom[ 2819]='h0000040c;  wr_data_rom[ 2819]='h00000000;
    rd_cycle[ 2820] = 1'b1;  wr_cycle[ 2820] = 1'b0;  addr_rom[ 2820]='h00000410;  wr_data_rom[ 2820]='h00000000;
    rd_cycle[ 2821] = 1'b1;  wr_cycle[ 2821] = 1'b0;  addr_rom[ 2821]='h00000414;  wr_data_rom[ 2821]='h00000000;
    rd_cycle[ 2822] = 1'b1;  wr_cycle[ 2822] = 1'b0;  addr_rom[ 2822]='h00000418;  wr_data_rom[ 2822]='h00000000;
    rd_cycle[ 2823] = 1'b1;  wr_cycle[ 2823] = 1'b0;  addr_rom[ 2823]='h0000041c;  wr_data_rom[ 2823]='h00000000;
    rd_cycle[ 2824] = 1'b1;  wr_cycle[ 2824] = 1'b0;  addr_rom[ 2824]='h00000420;  wr_data_rom[ 2824]='h00000000;
    rd_cycle[ 2825] = 1'b1;  wr_cycle[ 2825] = 1'b0;  addr_rom[ 2825]='h00000424;  wr_data_rom[ 2825]='h00000000;
    rd_cycle[ 2826] = 1'b1;  wr_cycle[ 2826] = 1'b0;  addr_rom[ 2826]='h00000428;  wr_data_rom[ 2826]='h00000000;
    rd_cycle[ 2827] = 1'b1;  wr_cycle[ 2827] = 1'b0;  addr_rom[ 2827]='h0000042c;  wr_data_rom[ 2827]='h00000000;
    rd_cycle[ 2828] = 1'b1;  wr_cycle[ 2828] = 1'b0;  addr_rom[ 2828]='h00000430;  wr_data_rom[ 2828]='h00000000;
    rd_cycle[ 2829] = 1'b1;  wr_cycle[ 2829] = 1'b0;  addr_rom[ 2829]='h00000434;  wr_data_rom[ 2829]='h00000000;
    rd_cycle[ 2830] = 1'b1;  wr_cycle[ 2830] = 1'b0;  addr_rom[ 2830]='h00000438;  wr_data_rom[ 2830]='h00000000;
    rd_cycle[ 2831] = 1'b1;  wr_cycle[ 2831] = 1'b0;  addr_rom[ 2831]='h0000043c;  wr_data_rom[ 2831]='h00000000;
    rd_cycle[ 2832] = 1'b1;  wr_cycle[ 2832] = 1'b0;  addr_rom[ 2832]='h00000440;  wr_data_rom[ 2832]='h00000000;
    rd_cycle[ 2833] = 1'b1;  wr_cycle[ 2833] = 1'b0;  addr_rom[ 2833]='h00000444;  wr_data_rom[ 2833]='h00000000;
    rd_cycle[ 2834] = 1'b1;  wr_cycle[ 2834] = 1'b0;  addr_rom[ 2834]='h00000448;  wr_data_rom[ 2834]='h00000000;
    rd_cycle[ 2835] = 1'b1;  wr_cycle[ 2835] = 1'b0;  addr_rom[ 2835]='h0000044c;  wr_data_rom[ 2835]='h00000000;
    rd_cycle[ 2836] = 1'b1;  wr_cycle[ 2836] = 1'b0;  addr_rom[ 2836]='h00000450;  wr_data_rom[ 2836]='h00000000;
    rd_cycle[ 2837] = 1'b1;  wr_cycle[ 2837] = 1'b0;  addr_rom[ 2837]='h00000454;  wr_data_rom[ 2837]='h00000000;
    rd_cycle[ 2838] = 1'b1;  wr_cycle[ 2838] = 1'b0;  addr_rom[ 2838]='h00000458;  wr_data_rom[ 2838]='h00000000;
    rd_cycle[ 2839] = 1'b1;  wr_cycle[ 2839] = 1'b0;  addr_rom[ 2839]='h0000045c;  wr_data_rom[ 2839]='h00000000;
    rd_cycle[ 2840] = 1'b1;  wr_cycle[ 2840] = 1'b0;  addr_rom[ 2840]='h00000460;  wr_data_rom[ 2840]='h00000000;
    rd_cycle[ 2841] = 1'b1;  wr_cycle[ 2841] = 1'b0;  addr_rom[ 2841]='h00000464;  wr_data_rom[ 2841]='h00000000;
    rd_cycle[ 2842] = 1'b1;  wr_cycle[ 2842] = 1'b0;  addr_rom[ 2842]='h00000468;  wr_data_rom[ 2842]='h00000000;
    rd_cycle[ 2843] = 1'b1;  wr_cycle[ 2843] = 1'b0;  addr_rom[ 2843]='h0000046c;  wr_data_rom[ 2843]='h00000000;
    rd_cycle[ 2844] = 1'b1;  wr_cycle[ 2844] = 1'b0;  addr_rom[ 2844]='h00000470;  wr_data_rom[ 2844]='h00000000;
    rd_cycle[ 2845] = 1'b1;  wr_cycle[ 2845] = 1'b0;  addr_rom[ 2845]='h00000474;  wr_data_rom[ 2845]='h00000000;
    rd_cycle[ 2846] = 1'b1;  wr_cycle[ 2846] = 1'b0;  addr_rom[ 2846]='h00000478;  wr_data_rom[ 2846]='h00000000;
    rd_cycle[ 2847] = 1'b1;  wr_cycle[ 2847] = 1'b0;  addr_rom[ 2847]='h0000047c;  wr_data_rom[ 2847]='h00000000;
    rd_cycle[ 2848] = 1'b1;  wr_cycle[ 2848] = 1'b0;  addr_rom[ 2848]='h00000480;  wr_data_rom[ 2848]='h00000000;
    rd_cycle[ 2849] = 1'b1;  wr_cycle[ 2849] = 1'b0;  addr_rom[ 2849]='h00000484;  wr_data_rom[ 2849]='h00000000;
    rd_cycle[ 2850] = 1'b1;  wr_cycle[ 2850] = 1'b0;  addr_rom[ 2850]='h00000488;  wr_data_rom[ 2850]='h00000000;
    rd_cycle[ 2851] = 1'b1;  wr_cycle[ 2851] = 1'b0;  addr_rom[ 2851]='h0000048c;  wr_data_rom[ 2851]='h00000000;
    rd_cycle[ 2852] = 1'b1;  wr_cycle[ 2852] = 1'b0;  addr_rom[ 2852]='h00000490;  wr_data_rom[ 2852]='h00000000;
    rd_cycle[ 2853] = 1'b1;  wr_cycle[ 2853] = 1'b0;  addr_rom[ 2853]='h00000494;  wr_data_rom[ 2853]='h00000000;
    rd_cycle[ 2854] = 1'b1;  wr_cycle[ 2854] = 1'b0;  addr_rom[ 2854]='h00000498;  wr_data_rom[ 2854]='h00000000;
    rd_cycle[ 2855] = 1'b1;  wr_cycle[ 2855] = 1'b0;  addr_rom[ 2855]='h0000049c;  wr_data_rom[ 2855]='h00000000;
    rd_cycle[ 2856] = 1'b1;  wr_cycle[ 2856] = 1'b0;  addr_rom[ 2856]='h000004a0;  wr_data_rom[ 2856]='h00000000;
    rd_cycle[ 2857] = 1'b1;  wr_cycle[ 2857] = 1'b0;  addr_rom[ 2857]='h000004a4;  wr_data_rom[ 2857]='h00000000;
    rd_cycle[ 2858] = 1'b1;  wr_cycle[ 2858] = 1'b0;  addr_rom[ 2858]='h000004a8;  wr_data_rom[ 2858]='h00000000;
    rd_cycle[ 2859] = 1'b1;  wr_cycle[ 2859] = 1'b0;  addr_rom[ 2859]='h000004ac;  wr_data_rom[ 2859]='h00000000;
    rd_cycle[ 2860] = 1'b1;  wr_cycle[ 2860] = 1'b0;  addr_rom[ 2860]='h000004b0;  wr_data_rom[ 2860]='h00000000;
    rd_cycle[ 2861] = 1'b1;  wr_cycle[ 2861] = 1'b0;  addr_rom[ 2861]='h000004b4;  wr_data_rom[ 2861]='h00000000;
    rd_cycle[ 2862] = 1'b1;  wr_cycle[ 2862] = 1'b0;  addr_rom[ 2862]='h000004b8;  wr_data_rom[ 2862]='h00000000;
    rd_cycle[ 2863] = 1'b1;  wr_cycle[ 2863] = 1'b0;  addr_rom[ 2863]='h000004bc;  wr_data_rom[ 2863]='h00000000;
    rd_cycle[ 2864] = 1'b1;  wr_cycle[ 2864] = 1'b0;  addr_rom[ 2864]='h000004c0;  wr_data_rom[ 2864]='h00000000;
    rd_cycle[ 2865] = 1'b1;  wr_cycle[ 2865] = 1'b0;  addr_rom[ 2865]='h000004c4;  wr_data_rom[ 2865]='h00000000;
    rd_cycle[ 2866] = 1'b1;  wr_cycle[ 2866] = 1'b0;  addr_rom[ 2866]='h000004c8;  wr_data_rom[ 2866]='h00000000;
    rd_cycle[ 2867] = 1'b1;  wr_cycle[ 2867] = 1'b0;  addr_rom[ 2867]='h000004cc;  wr_data_rom[ 2867]='h00000000;
    rd_cycle[ 2868] = 1'b1;  wr_cycle[ 2868] = 1'b0;  addr_rom[ 2868]='h000004d0;  wr_data_rom[ 2868]='h00000000;
    rd_cycle[ 2869] = 1'b1;  wr_cycle[ 2869] = 1'b0;  addr_rom[ 2869]='h000004d4;  wr_data_rom[ 2869]='h00000000;
    rd_cycle[ 2870] = 1'b1;  wr_cycle[ 2870] = 1'b0;  addr_rom[ 2870]='h000004d8;  wr_data_rom[ 2870]='h00000000;
    rd_cycle[ 2871] = 1'b1;  wr_cycle[ 2871] = 1'b0;  addr_rom[ 2871]='h000004dc;  wr_data_rom[ 2871]='h00000000;
    rd_cycle[ 2872] = 1'b1;  wr_cycle[ 2872] = 1'b0;  addr_rom[ 2872]='h000004e0;  wr_data_rom[ 2872]='h00000000;
    rd_cycle[ 2873] = 1'b1;  wr_cycle[ 2873] = 1'b0;  addr_rom[ 2873]='h000004e4;  wr_data_rom[ 2873]='h00000000;
    rd_cycle[ 2874] = 1'b1;  wr_cycle[ 2874] = 1'b0;  addr_rom[ 2874]='h000004e8;  wr_data_rom[ 2874]='h00000000;
    rd_cycle[ 2875] = 1'b1;  wr_cycle[ 2875] = 1'b0;  addr_rom[ 2875]='h000004ec;  wr_data_rom[ 2875]='h00000000;
    rd_cycle[ 2876] = 1'b1;  wr_cycle[ 2876] = 1'b0;  addr_rom[ 2876]='h000004f0;  wr_data_rom[ 2876]='h00000000;
    rd_cycle[ 2877] = 1'b1;  wr_cycle[ 2877] = 1'b0;  addr_rom[ 2877]='h000004f4;  wr_data_rom[ 2877]='h00000000;
    rd_cycle[ 2878] = 1'b1;  wr_cycle[ 2878] = 1'b0;  addr_rom[ 2878]='h000004f8;  wr_data_rom[ 2878]='h00000000;
    rd_cycle[ 2879] = 1'b1;  wr_cycle[ 2879] = 1'b0;  addr_rom[ 2879]='h000004fc;  wr_data_rom[ 2879]='h00000000;
    rd_cycle[ 2880] = 1'b1;  wr_cycle[ 2880] = 1'b0;  addr_rom[ 2880]='h00000500;  wr_data_rom[ 2880]='h00000000;
    rd_cycle[ 2881] = 1'b1;  wr_cycle[ 2881] = 1'b0;  addr_rom[ 2881]='h00000504;  wr_data_rom[ 2881]='h00000000;
    rd_cycle[ 2882] = 1'b1;  wr_cycle[ 2882] = 1'b0;  addr_rom[ 2882]='h00000508;  wr_data_rom[ 2882]='h00000000;
    rd_cycle[ 2883] = 1'b1;  wr_cycle[ 2883] = 1'b0;  addr_rom[ 2883]='h0000050c;  wr_data_rom[ 2883]='h00000000;
    rd_cycle[ 2884] = 1'b1;  wr_cycle[ 2884] = 1'b0;  addr_rom[ 2884]='h00000510;  wr_data_rom[ 2884]='h00000000;
    rd_cycle[ 2885] = 1'b1;  wr_cycle[ 2885] = 1'b0;  addr_rom[ 2885]='h00000514;  wr_data_rom[ 2885]='h00000000;
    rd_cycle[ 2886] = 1'b1;  wr_cycle[ 2886] = 1'b0;  addr_rom[ 2886]='h00000518;  wr_data_rom[ 2886]='h00000000;
    rd_cycle[ 2887] = 1'b1;  wr_cycle[ 2887] = 1'b0;  addr_rom[ 2887]='h0000051c;  wr_data_rom[ 2887]='h00000000;
    rd_cycle[ 2888] = 1'b1;  wr_cycle[ 2888] = 1'b0;  addr_rom[ 2888]='h00000520;  wr_data_rom[ 2888]='h00000000;
    rd_cycle[ 2889] = 1'b1;  wr_cycle[ 2889] = 1'b0;  addr_rom[ 2889]='h00000524;  wr_data_rom[ 2889]='h00000000;
    rd_cycle[ 2890] = 1'b1;  wr_cycle[ 2890] = 1'b0;  addr_rom[ 2890]='h00000528;  wr_data_rom[ 2890]='h00000000;
    rd_cycle[ 2891] = 1'b1;  wr_cycle[ 2891] = 1'b0;  addr_rom[ 2891]='h0000052c;  wr_data_rom[ 2891]='h00000000;
    rd_cycle[ 2892] = 1'b1;  wr_cycle[ 2892] = 1'b0;  addr_rom[ 2892]='h00000530;  wr_data_rom[ 2892]='h00000000;
    rd_cycle[ 2893] = 1'b1;  wr_cycle[ 2893] = 1'b0;  addr_rom[ 2893]='h00000534;  wr_data_rom[ 2893]='h00000000;
    rd_cycle[ 2894] = 1'b1;  wr_cycle[ 2894] = 1'b0;  addr_rom[ 2894]='h00000538;  wr_data_rom[ 2894]='h00000000;
    rd_cycle[ 2895] = 1'b1;  wr_cycle[ 2895] = 1'b0;  addr_rom[ 2895]='h0000053c;  wr_data_rom[ 2895]='h00000000;
    rd_cycle[ 2896] = 1'b1;  wr_cycle[ 2896] = 1'b0;  addr_rom[ 2896]='h00000540;  wr_data_rom[ 2896]='h00000000;
    rd_cycle[ 2897] = 1'b1;  wr_cycle[ 2897] = 1'b0;  addr_rom[ 2897]='h00000544;  wr_data_rom[ 2897]='h00000000;
    rd_cycle[ 2898] = 1'b1;  wr_cycle[ 2898] = 1'b0;  addr_rom[ 2898]='h00000548;  wr_data_rom[ 2898]='h00000000;
    rd_cycle[ 2899] = 1'b1;  wr_cycle[ 2899] = 1'b0;  addr_rom[ 2899]='h0000054c;  wr_data_rom[ 2899]='h00000000;
    rd_cycle[ 2900] = 1'b1;  wr_cycle[ 2900] = 1'b0;  addr_rom[ 2900]='h00000550;  wr_data_rom[ 2900]='h00000000;
    rd_cycle[ 2901] = 1'b1;  wr_cycle[ 2901] = 1'b0;  addr_rom[ 2901]='h00000554;  wr_data_rom[ 2901]='h00000000;
    rd_cycle[ 2902] = 1'b1;  wr_cycle[ 2902] = 1'b0;  addr_rom[ 2902]='h00000558;  wr_data_rom[ 2902]='h00000000;
    rd_cycle[ 2903] = 1'b1;  wr_cycle[ 2903] = 1'b0;  addr_rom[ 2903]='h0000055c;  wr_data_rom[ 2903]='h00000000;
    rd_cycle[ 2904] = 1'b1;  wr_cycle[ 2904] = 1'b0;  addr_rom[ 2904]='h00000560;  wr_data_rom[ 2904]='h00000000;
    rd_cycle[ 2905] = 1'b1;  wr_cycle[ 2905] = 1'b0;  addr_rom[ 2905]='h00000564;  wr_data_rom[ 2905]='h00000000;
    rd_cycle[ 2906] = 1'b1;  wr_cycle[ 2906] = 1'b0;  addr_rom[ 2906]='h00000568;  wr_data_rom[ 2906]='h00000000;
    rd_cycle[ 2907] = 1'b1;  wr_cycle[ 2907] = 1'b0;  addr_rom[ 2907]='h0000056c;  wr_data_rom[ 2907]='h00000000;
    rd_cycle[ 2908] = 1'b1;  wr_cycle[ 2908] = 1'b0;  addr_rom[ 2908]='h00000570;  wr_data_rom[ 2908]='h00000000;
    rd_cycle[ 2909] = 1'b1;  wr_cycle[ 2909] = 1'b0;  addr_rom[ 2909]='h00000574;  wr_data_rom[ 2909]='h00000000;
    rd_cycle[ 2910] = 1'b1;  wr_cycle[ 2910] = 1'b0;  addr_rom[ 2910]='h00000578;  wr_data_rom[ 2910]='h00000000;
    rd_cycle[ 2911] = 1'b1;  wr_cycle[ 2911] = 1'b0;  addr_rom[ 2911]='h0000057c;  wr_data_rom[ 2911]='h00000000;
    rd_cycle[ 2912] = 1'b1;  wr_cycle[ 2912] = 1'b0;  addr_rom[ 2912]='h00000580;  wr_data_rom[ 2912]='h00000000;
    rd_cycle[ 2913] = 1'b1;  wr_cycle[ 2913] = 1'b0;  addr_rom[ 2913]='h00000584;  wr_data_rom[ 2913]='h00000000;
    rd_cycle[ 2914] = 1'b1;  wr_cycle[ 2914] = 1'b0;  addr_rom[ 2914]='h00000588;  wr_data_rom[ 2914]='h00000000;
    rd_cycle[ 2915] = 1'b1;  wr_cycle[ 2915] = 1'b0;  addr_rom[ 2915]='h0000058c;  wr_data_rom[ 2915]='h00000000;
    rd_cycle[ 2916] = 1'b1;  wr_cycle[ 2916] = 1'b0;  addr_rom[ 2916]='h00000590;  wr_data_rom[ 2916]='h00000000;
    rd_cycle[ 2917] = 1'b1;  wr_cycle[ 2917] = 1'b0;  addr_rom[ 2917]='h00000594;  wr_data_rom[ 2917]='h00000000;
    rd_cycle[ 2918] = 1'b1;  wr_cycle[ 2918] = 1'b0;  addr_rom[ 2918]='h00000598;  wr_data_rom[ 2918]='h00000000;
    rd_cycle[ 2919] = 1'b1;  wr_cycle[ 2919] = 1'b0;  addr_rom[ 2919]='h0000059c;  wr_data_rom[ 2919]='h00000000;
    rd_cycle[ 2920] = 1'b1;  wr_cycle[ 2920] = 1'b0;  addr_rom[ 2920]='h000005a0;  wr_data_rom[ 2920]='h00000000;
    rd_cycle[ 2921] = 1'b1;  wr_cycle[ 2921] = 1'b0;  addr_rom[ 2921]='h000005a4;  wr_data_rom[ 2921]='h00000000;
    rd_cycle[ 2922] = 1'b1;  wr_cycle[ 2922] = 1'b0;  addr_rom[ 2922]='h000005a8;  wr_data_rom[ 2922]='h00000000;
    rd_cycle[ 2923] = 1'b1;  wr_cycle[ 2923] = 1'b0;  addr_rom[ 2923]='h000005ac;  wr_data_rom[ 2923]='h00000000;
    rd_cycle[ 2924] = 1'b1;  wr_cycle[ 2924] = 1'b0;  addr_rom[ 2924]='h000005b0;  wr_data_rom[ 2924]='h00000000;
    rd_cycle[ 2925] = 1'b1;  wr_cycle[ 2925] = 1'b0;  addr_rom[ 2925]='h000005b4;  wr_data_rom[ 2925]='h00000000;
    rd_cycle[ 2926] = 1'b1;  wr_cycle[ 2926] = 1'b0;  addr_rom[ 2926]='h000005b8;  wr_data_rom[ 2926]='h00000000;
    rd_cycle[ 2927] = 1'b1;  wr_cycle[ 2927] = 1'b0;  addr_rom[ 2927]='h000005bc;  wr_data_rom[ 2927]='h00000000;
    rd_cycle[ 2928] = 1'b1;  wr_cycle[ 2928] = 1'b0;  addr_rom[ 2928]='h000005c0;  wr_data_rom[ 2928]='h00000000;
    rd_cycle[ 2929] = 1'b1;  wr_cycle[ 2929] = 1'b0;  addr_rom[ 2929]='h000005c4;  wr_data_rom[ 2929]='h00000000;
    rd_cycle[ 2930] = 1'b1;  wr_cycle[ 2930] = 1'b0;  addr_rom[ 2930]='h000005c8;  wr_data_rom[ 2930]='h00000000;
    rd_cycle[ 2931] = 1'b1;  wr_cycle[ 2931] = 1'b0;  addr_rom[ 2931]='h000005cc;  wr_data_rom[ 2931]='h00000000;
    rd_cycle[ 2932] = 1'b1;  wr_cycle[ 2932] = 1'b0;  addr_rom[ 2932]='h000005d0;  wr_data_rom[ 2932]='h00000000;
    rd_cycle[ 2933] = 1'b1;  wr_cycle[ 2933] = 1'b0;  addr_rom[ 2933]='h000005d4;  wr_data_rom[ 2933]='h00000000;
    rd_cycle[ 2934] = 1'b1;  wr_cycle[ 2934] = 1'b0;  addr_rom[ 2934]='h000005d8;  wr_data_rom[ 2934]='h00000000;
    rd_cycle[ 2935] = 1'b1;  wr_cycle[ 2935] = 1'b0;  addr_rom[ 2935]='h000005dc;  wr_data_rom[ 2935]='h00000000;
    rd_cycle[ 2936] = 1'b1;  wr_cycle[ 2936] = 1'b0;  addr_rom[ 2936]='h000005e0;  wr_data_rom[ 2936]='h00000000;
    rd_cycle[ 2937] = 1'b1;  wr_cycle[ 2937] = 1'b0;  addr_rom[ 2937]='h000005e4;  wr_data_rom[ 2937]='h00000000;
    rd_cycle[ 2938] = 1'b1;  wr_cycle[ 2938] = 1'b0;  addr_rom[ 2938]='h000005e8;  wr_data_rom[ 2938]='h00000000;
    rd_cycle[ 2939] = 1'b1;  wr_cycle[ 2939] = 1'b0;  addr_rom[ 2939]='h000005ec;  wr_data_rom[ 2939]='h00000000;
    rd_cycle[ 2940] = 1'b1;  wr_cycle[ 2940] = 1'b0;  addr_rom[ 2940]='h000005f0;  wr_data_rom[ 2940]='h00000000;
    rd_cycle[ 2941] = 1'b1;  wr_cycle[ 2941] = 1'b0;  addr_rom[ 2941]='h000005f4;  wr_data_rom[ 2941]='h00000000;
    rd_cycle[ 2942] = 1'b1;  wr_cycle[ 2942] = 1'b0;  addr_rom[ 2942]='h000005f8;  wr_data_rom[ 2942]='h00000000;
    rd_cycle[ 2943] = 1'b1;  wr_cycle[ 2943] = 1'b0;  addr_rom[ 2943]='h000005fc;  wr_data_rom[ 2943]='h00000000;
    rd_cycle[ 2944] = 1'b1;  wr_cycle[ 2944] = 1'b0;  addr_rom[ 2944]='h00000600;  wr_data_rom[ 2944]='h00000000;
    rd_cycle[ 2945] = 1'b1;  wr_cycle[ 2945] = 1'b0;  addr_rom[ 2945]='h00000604;  wr_data_rom[ 2945]='h00000000;
    rd_cycle[ 2946] = 1'b1;  wr_cycle[ 2946] = 1'b0;  addr_rom[ 2946]='h00000608;  wr_data_rom[ 2946]='h00000000;
    rd_cycle[ 2947] = 1'b1;  wr_cycle[ 2947] = 1'b0;  addr_rom[ 2947]='h0000060c;  wr_data_rom[ 2947]='h00000000;
    rd_cycle[ 2948] = 1'b1;  wr_cycle[ 2948] = 1'b0;  addr_rom[ 2948]='h00000610;  wr_data_rom[ 2948]='h00000000;
    rd_cycle[ 2949] = 1'b1;  wr_cycle[ 2949] = 1'b0;  addr_rom[ 2949]='h00000614;  wr_data_rom[ 2949]='h00000000;
    rd_cycle[ 2950] = 1'b1;  wr_cycle[ 2950] = 1'b0;  addr_rom[ 2950]='h00000618;  wr_data_rom[ 2950]='h00000000;
    rd_cycle[ 2951] = 1'b1;  wr_cycle[ 2951] = 1'b0;  addr_rom[ 2951]='h0000061c;  wr_data_rom[ 2951]='h00000000;
    rd_cycle[ 2952] = 1'b1;  wr_cycle[ 2952] = 1'b0;  addr_rom[ 2952]='h00000620;  wr_data_rom[ 2952]='h00000000;
    rd_cycle[ 2953] = 1'b1;  wr_cycle[ 2953] = 1'b0;  addr_rom[ 2953]='h00000624;  wr_data_rom[ 2953]='h00000000;
    rd_cycle[ 2954] = 1'b1;  wr_cycle[ 2954] = 1'b0;  addr_rom[ 2954]='h00000628;  wr_data_rom[ 2954]='h00000000;
    rd_cycle[ 2955] = 1'b1;  wr_cycle[ 2955] = 1'b0;  addr_rom[ 2955]='h0000062c;  wr_data_rom[ 2955]='h00000000;
    rd_cycle[ 2956] = 1'b1;  wr_cycle[ 2956] = 1'b0;  addr_rom[ 2956]='h00000630;  wr_data_rom[ 2956]='h00000000;
    rd_cycle[ 2957] = 1'b1;  wr_cycle[ 2957] = 1'b0;  addr_rom[ 2957]='h00000634;  wr_data_rom[ 2957]='h00000000;
    rd_cycle[ 2958] = 1'b1;  wr_cycle[ 2958] = 1'b0;  addr_rom[ 2958]='h00000638;  wr_data_rom[ 2958]='h00000000;
    rd_cycle[ 2959] = 1'b1;  wr_cycle[ 2959] = 1'b0;  addr_rom[ 2959]='h0000063c;  wr_data_rom[ 2959]='h00000000;
    rd_cycle[ 2960] = 1'b1;  wr_cycle[ 2960] = 1'b0;  addr_rom[ 2960]='h00000640;  wr_data_rom[ 2960]='h00000000;
    rd_cycle[ 2961] = 1'b1;  wr_cycle[ 2961] = 1'b0;  addr_rom[ 2961]='h00000644;  wr_data_rom[ 2961]='h00000000;
    rd_cycle[ 2962] = 1'b1;  wr_cycle[ 2962] = 1'b0;  addr_rom[ 2962]='h00000648;  wr_data_rom[ 2962]='h00000000;
    rd_cycle[ 2963] = 1'b1;  wr_cycle[ 2963] = 1'b0;  addr_rom[ 2963]='h0000064c;  wr_data_rom[ 2963]='h00000000;
    rd_cycle[ 2964] = 1'b1;  wr_cycle[ 2964] = 1'b0;  addr_rom[ 2964]='h00000650;  wr_data_rom[ 2964]='h00000000;
    rd_cycle[ 2965] = 1'b1;  wr_cycle[ 2965] = 1'b0;  addr_rom[ 2965]='h00000654;  wr_data_rom[ 2965]='h00000000;
    rd_cycle[ 2966] = 1'b1;  wr_cycle[ 2966] = 1'b0;  addr_rom[ 2966]='h00000658;  wr_data_rom[ 2966]='h00000000;
    rd_cycle[ 2967] = 1'b1;  wr_cycle[ 2967] = 1'b0;  addr_rom[ 2967]='h0000065c;  wr_data_rom[ 2967]='h00000000;
    rd_cycle[ 2968] = 1'b1;  wr_cycle[ 2968] = 1'b0;  addr_rom[ 2968]='h00000660;  wr_data_rom[ 2968]='h00000000;
    rd_cycle[ 2969] = 1'b1;  wr_cycle[ 2969] = 1'b0;  addr_rom[ 2969]='h00000664;  wr_data_rom[ 2969]='h00000000;
    rd_cycle[ 2970] = 1'b1;  wr_cycle[ 2970] = 1'b0;  addr_rom[ 2970]='h00000668;  wr_data_rom[ 2970]='h00000000;
    rd_cycle[ 2971] = 1'b1;  wr_cycle[ 2971] = 1'b0;  addr_rom[ 2971]='h0000066c;  wr_data_rom[ 2971]='h00000000;
    rd_cycle[ 2972] = 1'b1;  wr_cycle[ 2972] = 1'b0;  addr_rom[ 2972]='h00000670;  wr_data_rom[ 2972]='h00000000;
    rd_cycle[ 2973] = 1'b1;  wr_cycle[ 2973] = 1'b0;  addr_rom[ 2973]='h00000674;  wr_data_rom[ 2973]='h00000000;
    rd_cycle[ 2974] = 1'b1;  wr_cycle[ 2974] = 1'b0;  addr_rom[ 2974]='h00000678;  wr_data_rom[ 2974]='h00000000;
    rd_cycle[ 2975] = 1'b1;  wr_cycle[ 2975] = 1'b0;  addr_rom[ 2975]='h0000067c;  wr_data_rom[ 2975]='h00000000;
    rd_cycle[ 2976] = 1'b1;  wr_cycle[ 2976] = 1'b0;  addr_rom[ 2976]='h00000680;  wr_data_rom[ 2976]='h00000000;
    rd_cycle[ 2977] = 1'b1;  wr_cycle[ 2977] = 1'b0;  addr_rom[ 2977]='h00000684;  wr_data_rom[ 2977]='h00000000;
    rd_cycle[ 2978] = 1'b1;  wr_cycle[ 2978] = 1'b0;  addr_rom[ 2978]='h00000688;  wr_data_rom[ 2978]='h00000000;
    rd_cycle[ 2979] = 1'b1;  wr_cycle[ 2979] = 1'b0;  addr_rom[ 2979]='h0000068c;  wr_data_rom[ 2979]='h00000000;
    rd_cycle[ 2980] = 1'b1;  wr_cycle[ 2980] = 1'b0;  addr_rom[ 2980]='h00000690;  wr_data_rom[ 2980]='h00000000;
    rd_cycle[ 2981] = 1'b1;  wr_cycle[ 2981] = 1'b0;  addr_rom[ 2981]='h00000694;  wr_data_rom[ 2981]='h00000000;
    rd_cycle[ 2982] = 1'b1;  wr_cycle[ 2982] = 1'b0;  addr_rom[ 2982]='h00000698;  wr_data_rom[ 2982]='h00000000;
    rd_cycle[ 2983] = 1'b1;  wr_cycle[ 2983] = 1'b0;  addr_rom[ 2983]='h0000069c;  wr_data_rom[ 2983]='h00000000;
    rd_cycle[ 2984] = 1'b1;  wr_cycle[ 2984] = 1'b0;  addr_rom[ 2984]='h000006a0;  wr_data_rom[ 2984]='h00000000;
    rd_cycle[ 2985] = 1'b1;  wr_cycle[ 2985] = 1'b0;  addr_rom[ 2985]='h000006a4;  wr_data_rom[ 2985]='h00000000;
    rd_cycle[ 2986] = 1'b1;  wr_cycle[ 2986] = 1'b0;  addr_rom[ 2986]='h000006a8;  wr_data_rom[ 2986]='h00000000;
    rd_cycle[ 2987] = 1'b1;  wr_cycle[ 2987] = 1'b0;  addr_rom[ 2987]='h000006ac;  wr_data_rom[ 2987]='h00000000;
    rd_cycle[ 2988] = 1'b1;  wr_cycle[ 2988] = 1'b0;  addr_rom[ 2988]='h000006b0;  wr_data_rom[ 2988]='h00000000;
    rd_cycle[ 2989] = 1'b1;  wr_cycle[ 2989] = 1'b0;  addr_rom[ 2989]='h000006b4;  wr_data_rom[ 2989]='h00000000;
    rd_cycle[ 2990] = 1'b1;  wr_cycle[ 2990] = 1'b0;  addr_rom[ 2990]='h000006b8;  wr_data_rom[ 2990]='h00000000;
    rd_cycle[ 2991] = 1'b1;  wr_cycle[ 2991] = 1'b0;  addr_rom[ 2991]='h000006bc;  wr_data_rom[ 2991]='h00000000;
    rd_cycle[ 2992] = 1'b1;  wr_cycle[ 2992] = 1'b0;  addr_rom[ 2992]='h000006c0;  wr_data_rom[ 2992]='h00000000;
    rd_cycle[ 2993] = 1'b1;  wr_cycle[ 2993] = 1'b0;  addr_rom[ 2993]='h000006c4;  wr_data_rom[ 2993]='h00000000;
    rd_cycle[ 2994] = 1'b1;  wr_cycle[ 2994] = 1'b0;  addr_rom[ 2994]='h000006c8;  wr_data_rom[ 2994]='h00000000;
    rd_cycle[ 2995] = 1'b1;  wr_cycle[ 2995] = 1'b0;  addr_rom[ 2995]='h000006cc;  wr_data_rom[ 2995]='h00000000;
    rd_cycle[ 2996] = 1'b1;  wr_cycle[ 2996] = 1'b0;  addr_rom[ 2996]='h000006d0;  wr_data_rom[ 2996]='h00000000;
    rd_cycle[ 2997] = 1'b1;  wr_cycle[ 2997] = 1'b0;  addr_rom[ 2997]='h000006d4;  wr_data_rom[ 2997]='h00000000;
    rd_cycle[ 2998] = 1'b1;  wr_cycle[ 2998] = 1'b0;  addr_rom[ 2998]='h000006d8;  wr_data_rom[ 2998]='h00000000;
    rd_cycle[ 2999] = 1'b1;  wr_cycle[ 2999] = 1'b0;  addr_rom[ 2999]='h000006dc;  wr_data_rom[ 2999]='h00000000;
    rd_cycle[ 3000] = 1'b1;  wr_cycle[ 3000] = 1'b0;  addr_rom[ 3000]='h000006e0;  wr_data_rom[ 3000]='h00000000;
    rd_cycle[ 3001] = 1'b1;  wr_cycle[ 3001] = 1'b0;  addr_rom[ 3001]='h000006e4;  wr_data_rom[ 3001]='h00000000;
    rd_cycle[ 3002] = 1'b1;  wr_cycle[ 3002] = 1'b0;  addr_rom[ 3002]='h000006e8;  wr_data_rom[ 3002]='h00000000;
    rd_cycle[ 3003] = 1'b1;  wr_cycle[ 3003] = 1'b0;  addr_rom[ 3003]='h000006ec;  wr_data_rom[ 3003]='h00000000;
    rd_cycle[ 3004] = 1'b1;  wr_cycle[ 3004] = 1'b0;  addr_rom[ 3004]='h000006f0;  wr_data_rom[ 3004]='h00000000;
    rd_cycle[ 3005] = 1'b1;  wr_cycle[ 3005] = 1'b0;  addr_rom[ 3005]='h000006f4;  wr_data_rom[ 3005]='h00000000;
    rd_cycle[ 3006] = 1'b1;  wr_cycle[ 3006] = 1'b0;  addr_rom[ 3006]='h000006f8;  wr_data_rom[ 3006]='h00000000;
    rd_cycle[ 3007] = 1'b1;  wr_cycle[ 3007] = 1'b0;  addr_rom[ 3007]='h000006fc;  wr_data_rom[ 3007]='h00000000;
    rd_cycle[ 3008] = 1'b1;  wr_cycle[ 3008] = 1'b0;  addr_rom[ 3008]='h00000700;  wr_data_rom[ 3008]='h00000000;
    rd_cycle[ 3009] = 1'b1;  wr_cycle[ 3009] = 1'b0;  addr_rom[ 3009]='h00000704;  wr_data_rom[ 3009]='h00000000;
    rd_cycle[ 3010] = 1'b1;  wr_cycle[ 3010] = 1'b0;  addr_rom[ 3010]='h00000708;  wr_data_rom[ 3010]='h00000000;
    rd_cycle[ 3011] = 1'b1;  wr_cycle[ 3011] = 1'b0;  addr_rom[ 3011]='h0000070c;  wr_data_rom[ 3011]='h00000000;
    rd_cycle[ 3012] = 1'b1;  wr_cycle[ 3012] = 1'b0;  addr_rom[ 3012]='h00000710;  wr_data_rom[ 3012]='h00000000;
    rd_cycle[ 3013] = 1'b1;  wr_cycle[ 3013] = 1'b0;  addr_rom[ 3013]='h00000714;  wr_data_rom[ 3013]='h00000000;
    rd_cycle[ 3014] = 1'b1;  wr_cycle[ 3014] = 1'b0;  addr_rom[ 3014]='h00000718;  wr_data_rom[ 3014]='h00000000;
    rd_cycle[ 3015] = 1'b1;  wr_cycle[ 3015] = 1'b0;  addr_rom[ 3015]='h0000071c;  wr_data_rom[ 3015]='h00000000;
    rd_cycle[ 3016] = 1'b1;  wr_cycle[ 3016] = 1'b0;  addr_rom[ 3016]='h00000720;  wr_data_rom[ 3016]='h00000000;
    rd_cycle[ 3017] = 1'b1;  wr_cycle[ 3017] = 1'b0;  addr_rom[ 3017]='h00000724;  wr_data_rom[ 3017]='h00000000;
    rd_cycle[ 3018] = 1'b1;  wr_cycle[ 3018] = 1'b0;  addr_rom[ 3018]='h00000728;  wr_data_rom[ 3018]='h00000000;
    rd_cycle[ 3019] = 1'b1;  wr_cycle[ 3019] = 1'b0;  addr_rom[ 3019]='h0000072c;  wr_data_rom[ 3019]='h00000000;
    rd_cycle[ 3020] = 1'b1;  wr_cycle[ 3020] = 1'b0;  addr_rom[ 3020]='h00000730;  wr_data_rom[ 3020]='h00000000;
    rd_cycle[ 3021] = 1'b1;  wr_cycle[ 3021] = 1'b0;  addr_rom[ 3021]='h00000734;  wr_data_rom[ 3021]='h00000000;
    rd_cycle[ 3022] = 1'b1;  wr_cycle[ 3022] = 1'b0;  addr_rom[ 3022]='h00000738;  wr_data_rom[ 3022]='h00000000;
    rd_cycle[ 3023] = 1'b1;  wr_cycle[ 3023] = 1'b0;  addr_rom[ 3023]='h0000073c;  wr_data_rom[ 3023]='h00000000;
    rd_cycle[ 3024] = 1'b1;  wr_cycle[ 3024] = 1'b0;  addr_rom[ 3024]='h00000740;  wr_data_rom[ 3024]='h00000000;
    rd_cycle[ 3025] = 1'b1;  wr_cycle[ 3025] = 1'b0;  addr_rom[ 3025]='h00000744;  wr_data_rom[ 3025]='h00000000;
    rd_cycle[ 3026] = 1'b1;  wr_cycle[ 3026] = 1'b0;  addr_rom[ 3026]='h00000748;  wr_data_rom[ 3026]='h00000000;
    rd_cycle[ 3027] = 1'b1;  wr_cycle[ 3027] = 1'b0;  addr_rom[ 3027]='h0000074c;  wr_data_rom[ 3027]='h00000000;
    rd_cycle[ 3028] = 1'b1;  wr_cycle[ 3028] = 1'b0;  addr_rom[ 3028]='h00000750;  wr_data_rom[ 3028]='h00000000;
    rd_cycle[ 3029] = 1'b1;  wr_cycle[ 3029] = 1'b0;  addr_rom[ 3029]='h00000754;  wr_data_rom[ 3029]='h00000000;
    rd_cycle[ 3030] = 1'b1;  wr_cycle[ 3030] = 1'b0;  addr_rom[ 3030]='h00000758;  wr_data_rom[ 3030]='h00000000;
    rd_cycle[ 3031] = 1'b1;  wr_cycle[ 3031] = 1'b0;  addr_rom[ 3031]='h0000075c;  wr_data_rom[ 3031]='h00000000;
    rd_cycle[ 3032] = 1'b1;  wr_cycle[ 3032] = 1'b0;  addr_rom[ 3032]='h00000760;  wr_data_rom[ 3032]='h00000000;
    rd_cycle[ 3033] = 1'b1;  wr_cycle[ 3033] = 1'b0;  addr_rom[ 3033]='h00000764;  wr_data_rom[ 3033]='h00000000;
    rd_cycle[ 3034] = 1'b1;  wr_cycle[ 3034] = 1'b0;  addr_rom[ 3034]='h00000768;  wr_data_rom[ 3034]='h00000000;
    rd_cycle[ 3035] = 1'b1;  wr_cycle[ 3035] = 1'b0;  addr_rom[ 3035]='h0000076c;  wr_data_rom[ 3035]='h00000000;
    rd_cycle[ 3036] = 1'b1;  wr_cycle[ 3036] = 1'b0;  addr_rom[ 3036]='h00000770;  wr_data_rom[ 3036]='h00000000;
    rd_cycle[ 3037] = 1'b1;  wr_cycle[ 3037] = 1'b0;  addr_rom[ 3037]='h00000774;  wr_data_rom[ 3037]='h00000000;
    rd_cycle[ 3038] = 1'b1;  wr_cycle[ 3038] = 1'b0;  addr_rom[ 3038]='h00000778;  wr_data_rom[ 3038]='h00000000;
    rd_cycle[ 3039] = 1'b1;  wr_cycle[ 3039] = 1'b0;  addr_rom[ 3039]='h0000077c;  wr_data_rom[ 3039]='h00000000;
    rd_cycle[ 3040] = 1'b1;  wr_cycle[ 3040] = 1'b0;  addr_rom[ 3040]='h00000780;  wr_data_rom[ 3040]='h00000000;
    rd_cycle[ 3041] = 1'b1;  wr_cycle[ 3041] = 1'b0;  addr_rom[ 3041]='h00000784;  wr_data_rom[ 3041]='h00000000;
    rd_cycle[ 3042] = 1'b1;  wr_cycle[ 3042] = 1'b0;  addr_rom[ 3042]='h00000788;  wr_data_rom[ 3042]='h00000000;
    rd_cycle[ 3043] = 1'b1;  wr_cycle[ 3043] = 1'b0;  addr_rom[ 3043]='h0000078c;  wr_data_rom[ 3043]='h00000000;
    rd_cycle[ 3044] = 1'b1;  wr_cycle[ 3044] = 1'b0;  addr_rom[ 3044]='h00000790;  wr_data_rom[ 3044]='h00000000;
    rd_cycle[ 3045] = 1'b1;  wr_cycle[ 3045] = 1'b0;  addr_rom[ 3045]='h00000794;  wr_data_rom[ 3045]='h00000000;
    rd_cycle[ 3046] = 1'b1;  wr_cycle[ 3046] = 1'b0;  addr_rom[ 3046]='h00000798;  wr_data_rom[ 3046]='h00000000;
    rd_cycle[ 3047] = 1'b1;  wr_cycle[ 3047] = 1'b0;  addr_rom[ 3047]='h0000079c;  wr_data_rom[ 3047]='h00000000;
    rd_cycle[ 3048] = 1'b1;  wr_cycle[ 3048] = 1'b0;  addr_rom[ 3048]='h000007a0;  wr_data_rom[ 3048]='h00000000;
    rd_cycle[ 3049] = 1'b1;  wr_cycle[ 3049] = 1'b0;  addr_rom[ 3049]='h000007a4;  wr_data_rom[ 3049]='h00000000;
    rd_cycle[ 3050] = 1'b1;  wr_cycle[ 3050] = 1'b0;  addr_rom[ 3050]='h000007a8;  wr_data_rom[ 3050]='h00000000;
    rd_cycle[ 3051] = 1'b1;  wr_cycle[ 3051] = 1'b0;  addr_rom[ 3051]='h000007ac;  wr_data_rom[ 3051]='h00000000;
    rd_cycle[ 3052] = 1'b1;  wr_cycle[ 3052] = 1'b0;  addr_rom[ 3052]='h000007b0;  wr_data_rom[ 3052]='h00000000;
    rd_cycle[ 3053] = 1'b1;  wr_cycle[ 3053] = 1'b0;  addr_rom[ 3053]='h000007b4;  wr_data_rom[ 3053]='h00000000;
    rd_cycle[ 3054] = 1'b1;  wr_cycle[ 3054] = 1'b0;  addr_rom[ 3054]='h000007b8;  wr_data_rom[ 3054]='h00000000;
    rd_cycle[ 3055] = 1'b1;  wr_cycle[ 3055] = 1'b0;  addr_rom[ 3055]='h000007bc;  wr_data_rom[ 3055]='h00000000;
    rd_cycle[ 3056] = 1'b1;  wr_cycle[ 3056] = 1'b0;  addr_rom[ 3056]='h000007c0;  wr_data_rom[ 3056]='h00000000;
    rd_cycle[ 3057] = 1'b1;  wr_cycle[ 3057] = 1'b0;  addr_rom[ 3057]='h000007c4;  wr_data_rom[ 3057]='h00000000;
    rd_cycle[ 3058] = 1'b1;  wr_cycle[ 3058] = 1'b0;  addr_rom[ 3058]='h000007c8;  wr_data_rom[ 3058]='h00000000;
    rd_cycle[ 3059] = 1'b1;  wr_cycle[ 3059] = 1'b0;  addr_rom[ 3059]='h000007cc;  wr_data_rom[ 3059]='h00000000;
    rd_cycle[ 3060] = 1'b1;  wr_cycle[ 3060] = 1'b0;  addr_rom[ 3060]='h000007d0;  wr_data_rom[ 3060]='h00000000;
    rd_cycle[ 3061] = 1'b1;  wr_cycle[ 3061] = 1'b0;  addr_rom[ 3061]='h000007d4;  wr_data_rom[ 3061]='h00000000;
    rd_cycle[ 3062] = 1'b1;  wr_cycle[ 3062] = 1'b0;  addr_rom[ 3062]='h000007d8;  wr_data_rom[ 3062]='h00000000;
    rd_cycle[ 3063] = 1'b1;  wr_cycle[ 3063] = 1'b0;  addr_rom[ 3063]='h000007dc;  wr_data_rom[ 3063]='h00000000;
    rd_cycle[ 3064] = 1'b1;  wr_cycle[ 3064] = 1'b0;  addr_rom[ 3064]='h000007e0;  wr_data_rom[ 3064]='h00000000;
    rd_cycle[ 3065] = 1'b1;  wr_cycle[ 3065] = 1'b0;  addr_rom[ 3065]='h000007e4;  wr_data_rom[ 3065]='h00000000;
    rd_cycle[ 3066] = 1'b1;  wr_cycle[ 3066] = 1'b0;  addr_rom[ 3066]='h000007e8;  wr_data_rom[ 3066]='h00000000;
    rd_cycle[ 3067] = 1'b1;  wr_cycle[ 3067] = 1'b0;  addr_rom[ 3067]='h000007ec;  wr_data_rom[ 3067]='h00000000;
    rd_cycle[ 3068] = 1'b1;  wr_cycle[ 3068] = 1'b0;  addr_rom[ 3068]='h000007f0;  wr_data_rom[ 3068]='h00000000;
    rd_cycle[ 3069] = 1'b1;  wr_cycle[ 3069] = 1'b0;  addr_rom[ 3069]='h000007f4;  wr_data_rom[ 3069]='h00000000;
    rd_cycle[ 3070] = 1'b1;  wr_cycle[ 3070] = 1'b0;  addr_rom[ 3070]='h000007f8;  wr_data_rom[ 3070]='h00000000;
    rd_cycle[ 3071] = 1'b1;  wr_cycle[ 3071] = 1'b0;  addr_rom[ 3071]='h000007fc;  wr_data_rom[ 3071]='h00000000;
end

initial begin
    validation_data[    0] = 'h000004dd; 
    validation_data[    1] = 'h000006c4; 
    validation_data[    2] = 'h000006de; 
    validation_data[    3] = 'h000003bb; 
    validation_data[    4] = 'h000006db; 
    validation_data[    5] = 'h000006d7; 
    validation_data[    6] = 'h0000027c; 
    validation_data[    7] = 'h00000278; 
    validation_data[    8] = 'h00000628; 
    validation_data[    9] = 'h00000646; 
    validation_data[   10] = 'h00000590; 
    validation_data[   11] = 'h0000039d; 
    validation_data[   12] = 'h00000472; 
    validation_data[   13] = 'h00000780; 
    validation_data[   14] = 'h000001a3; 
    validation_data[   15] = 'h00000031; 
    validation_data[   16] = 'h0000000e; 
    validation_data[   17] = 'h00000266; 
    validation_data[   18] = 'h00000578; 
    validation_data[   19] = 'h000003e1; 
    validation_data[   20] = 'h000003c4; 
    validation_data[   21] = 'h00000377; 
    validation_data[   22] = 'h00000288; 
    validation_data[   23] = 'h000001e2; 
    validation_data[   24] = 'h00000224; 
    validation_data[   25] = 'h000001da; 
    validation_data[   26] = 'h00000765; 
    validation_data[   27] = 'h000006c4; 
    validation_data[   28] = 'h0000036b; 
    validation_data[   29] = 'h00000753; 
    validation_data[   30] = 'h00000058; 
    validation_data[   31] = 'h00000526; 
    validation_data[   32] = 'h000004be; 
    validation_data[   33] = 'h000003a5; 
    validation_data[   34] = 'h0000045a; 
    validation_data[   35] = 'h000003bb; 
    validation_data[   36] = 'h0000068a; 
    validation_data[   37] = 'h00000547; 
    validation_data[   38] = 'h000002af; 
    validation_data[   39] = 'h00000533; 
    validation_data[   40] = 'h000000af; 
    validation_data[   41] = 'h00000290; 
    validation_data[   42] = 'h00000688; 
    validation_data[   43] = 'h00000654; 
    validation_data[   44] = 'h00000771; 
    validation_data[   45] = 'h0000011a; 
    validation_data[   46] = 'h00000012; 
    validation_data[   47] = 'h000007c2; 
    validation_data[   48] = 'h0000007c; 
    validation_data[   49] = 'h000000b5; 
    validation_data[   50] = 'h0000011f; 
    validation_data[   51] = 'h000003d8; 
    validation_data[   52] = 'h0000061a; 
    validation_data[   53] = 'h000003d0; 
    validation_data[   54] = 'h000000c2; 
    validation_data[   55] = 'h000002af; 
    validation_data[   56] = 'h0000055f; 
    validation_data[   57] = 'h00000763; 
    validation_data[   58] = 'h000001aa; 
    validation_data[   59] = 'h000003d7; 
    validation_data[   60] = 'h000000be; 
    validation_data[   61] = 'h00000767; 
    validation_data[   62] = 'h000007e9; 
    validation_data[   63] = 'h00000741; 
    validation_data[   64] = 'h000000a9; 
    validation_data[   65] = 'h0000069a; 
    validation_data[   66] = 'h00000406; 
    validation_data[   67] = 'h00000083; 
    validation_data[   68] = 'h0000012f; 
    validation_data[   69] = 'h00000316; 
    validation_data[   70] = 'h000004a9; 
    validation_data[   71] = 'h000006b1; 
    validation_data[   72] = 'h000002bb; 
    validation_data[   73] = 'h000001fb; 
    validation_data[   74] = 'h0000053f; 
    validation_data[   75] = 'h0000033b; 
    validation_data[   76] = 'h00000002; 
    validation_data[   77] = 'h0000011d; 
    validation_data[   78] = 'h0000061a; 
    validation_data[   79] = 'h0000005d; 
    validation_data[   80] = 'h000003fc; 
    validation_data[   81] = 'h000004a6; 
    validation_data[   82] = 'h000001cb; 
    validation_data[   83] = 'h00000273; 
    validation_data[   84] = 'h000003b1; 
    validation_data[   85] = 'h00000084; 
    validation_data[   86] = 'h000000e2; 
    validation_data[   87] = 'h00000089; 
    validation_data[   88] = 'h00000519; 
    validation_data[   89] = 'h0000044e; 
    validation_data[   90] = 'h000004cf; 
    validation_data[   91] = 'h000001f5; 
    validation_data[   92] = 'h000004c0; 
    validation_data[   93] = 'h00000312; 
    validation_data[   94] = 'h00000049; 
    validation_data[   95] = 'h000002ba; 
    validation_data[   96] = 'h0000074e; 
    validation_data[   97] = 'h00000390; 
    validation_data[   98] = 'h0000065e; 
    validation_data[   99] = 'h000000c8; 
    validation_data[  100] = 'h0000008e; 
    validation_data[  101] = 'h0000015b; 
    validation_data[  102] = 'h000006a7; 
    validation_data[  103] = 'h000000da; 
    validation_data[  104] = 'h0000029d; 
    validation_data[  105] = 'h00000281; 
    validation_data[  106] = 'h000004eb; 
    validation_data[  107] = 'h00000704; 
    validation_data[  108] = 'h000007aa; 
    validation_data[  109] = 'h0000022e; 
    validation_data[  110] = 'h000004c5; 
    validation_data[  111] = 'h00000241; 
    validation_data[  112] = 'h00000071; 
    validation_data[  113] = 'h000003b4; 
    validation_data[  114] = 'h00000534; 
    validation_data[  115] = 'h0000042d; 
    validation_data[  116] = 'h000000a0; 
    validation_data[  117] = 'h00000488; 
    validation_data[  118] = 'h000000f2; 
    validation_data[  119] = 'h00000170; 
    validation_data[  120] = 'h00000441; 
    validation_data[  121] = 'h0000004d; 
    validation_data[  122] = 'h00000514; 
    validation_data[  123] = 'h00000781; 
    validation_data[  124] = 'h000007f0; 
    validation_data[  125] = 'h0000074b; 
    validation_data[  126] = 'h000004eb; 
    validation_data[  127] = 'h0000024f; 
    validation_data[  128] = 'h000002c9; 
    validation_data[  129] = 'h000002c1; 
    validation_data[  130] = 'h0000028e; 
    validation_data[  131] = 'h00000549; 
    validation_data[  132] = 'h000001af; 
    validation_data[  133] = 'h000001d5; 
    validation_data[  134] = 'h000003ad; 
    validation_data[  135] = 'h00000635; 
    validation_data[  136] = 'h0000018c; 
    validation_data[  137] = 'h000006e5; 
    validation_data[  138] = 'h00000432; 
    validation_data[  139] = 'h00000530; 
    validation_data[  140] = 'h0000019e; 
    validation_data[  141] = 'h00000588; 
    validation_data[  142] = 'h000003c9; 
    validation_data[  143] = 'h0000043d; 
    validation_data[  144] = 'h0000061e; 
    validation_data[  145] = 'h0000023a; 
    validation_data[  146] = 'h000000aa; 
    validation_data[  147] = 'h00000203; 
    validation_data[  148] = 'h0000056f; 
    validation_data[  149] = 'h000004b5; 
    validation_data[  150] = 'h000002b2; 
    validation_data[  151] = 'h000002e3; 
    validation_data[  152] = 'h000007d9; 
    validation_data[  153] = 'h000001c6; 
    validation_data[  154] = 'h00000290; 
    validation_data[  155] = 'h000002e7; 
    validation_data[  156] = 'h000001f9; 
    validation_data[  157] = 'h000001dd; 
    validation_data[  158] = 'h00000041; 
    validation_data[  159] = 'h000001e1; 
    validation_data[  160] = 'h00000402; 
    validation_data[  161] = 'h000002bd; 
    validation_data[  162] = 'h000004b9; 
    validation_data[  163] = 'h00000595; 
    validation_data[  164] = 'h00000740; 
    validation_data[  165] = 'h000002be; 
    validation_data[  166] = 'h00000699; 
    validation_data[  167] = 'h0000073d; 
    validation_data[  168] = 'h0000020d; 
    validation_data[  169] = 'h0000024b; 
    validation_data[  170] = 'h0000059e; 
    validation_data[  171] = 'h0000035f; 
    validation_data[  172] = 'h00000241; 
    validation_data[  173] = 'h00000288; 
    validation_data[  174] = 'h00000479; 
    validation_data[  175] = 'h000002b4; 
    validation_data[  176] = 'h000000a9; 
    validation_data[  177] = 'h00000555; 
    validation_data[  178] = 'h000002f7; 
    validation_data[  179] = 'h0000003b; 
    validation_data[  180] = 'h0000067b; 
    validation_data[  181] = 'h000002b4; 
    validation_data[  182] = 'h00000327; 
    validation_data[  183] = 'h0000012a; 
    validation_data[  184] = 'h000001a6; 
    validation_data[  185] = 'h000005cf; 
    validation_data[  186] = 'h000000da; 
    validation_data[  187] = 'h0000025d; 
    validation_data[  188] = 'h0000018d; 
    validation_data[  189] = 'h000003c5; 
    validation_data[  190] = 'h0000078b; 
    validation_data[  191] = 'h00000215; 
    validation_data[  192] = 'h0000033e; 
    validation_data[  193] = 'h0000068a; 
    validation_data[  194] = 'h0000076c; 
    validation_data[  195] = 'h00000712; 
    validation_data[  196] = 'h00000589; 
    validation_data[  197] = 'h00000778; 
    validation_data[  198] = 'h000003fa; 
    validation_data[  199] = 'h00000546; 
    validation_data[  200] = 'h000002d9; 
    validation_data[  201] = 'h000005e8; 
    validation_data[  202] = 'h0000059d; 
    validation_data[  203] = 'h00000235; 
    validation_data[  204] = 'h000003cb; 
    validation_data[  205] = 'h000002ba; 
    validation_data[  206] = 'h00000670; 
    validation_data[  207] = 'h00000150; 
    validation_data[  208] = 'h0000077a; 
    validation_data[  209] = 'h00000530; 
    validation_data[  210] = 'h0000070a; 
    validation_data[  211] = 'h00000143; 
    validation_data[  212] = 'h000006e7; 
    validation_data[  213] = 'h00000116; 
    validation_data[  214] = 'h0000031d; 
    validation_data[  215] = 'h000007e1; 
    validation_data[  216] = 'h000005dd; 
    validation_data[  217] = 'h00000031; 
    validation_data[  218] = 'h000003bf; 
    validation_data[  219] = 'h0000051a; 
    validation_data[  220] = 'h000006e8; 
    validation_data[  221] = 'h00000244; 
    validation_data[  222] = 'h000000a5; 
    validation_data[  223] = 'h000005e4; 
    validation_data[  224] = 'h00000597; 
    validation_data[  225] = 'h000004c0; 
    validation_data[  226] = 'h000006cb; 
    validation_data[  227] = 'h000007ca; 
    validation_data[  228] = 'h0000014f; 
    validation_data[  229] = 'h00000555; 
    validation_data[  230] = 'h000003d0; 
    validation_data[  231] = 'h00000374; 
    validation_data[  232] = 'h0000046a; 
    validation_data[  233] = 'h00000344; 
    validation_data[  234] = 'h00000111; 
    validation_data[  235] = 'h00000210; 
    validation_data[  236] = 'h000007a3; 
    validation_data[  237] = 'h0000001d; 
    validation_data[  238] = 'h00000587; 
    validation_data[  239] = 'h000002a5; 
    validation_data[  240] = 'h0000042a; 
    validation_data[  241] = 'h000000d6; 
    validation_data[  242] = 'h000003d3; 
    validation_data[  243] = 'h0000072e; 
    validation_data[  244] = 'h000004d6; 
    validation_data[  245] = 'h0000001e; 
    validation_data[  246] = 'h00000677; 
    validation_data[  247] = 'h0000007b; 
    validation_data[  248] = 'h0000044a; 
    validation_data[  249] = 'h000007d1; 
    validation_data[  250] = 'h00000224; 
    validation_data[  251] = 'h00000210; 
    validation_data[  252] = 'h0000011f; 
    validation_data[  253] = 'h000005ed; 
    validation_data[  254] = 'h00000243; 
    validation_data[  255] = 'h00000223; 
    validation_data[  256] = 'h00000382; 
    validation_data[  257] = 'h00000453; 
    validation_data[  258] = 'h00000050; 
    validation_data[  259] = 'h000001db; 
    validation_data[  260] = 'h00000227; 
    validation_data[  261] = 'h000001c2; 
    validation_data[  262] = 'h000005df; 
    validation_data[  263] = 'h000002ac; 
    validation_data[  264] = 'h00000595; 
    validation_data[  265] = 'h00000057; 
    validation_data[  266] = 'h0000029a; 
    validation_data[  267] = 'h000003f7; 
    validation_data[  268] = 'h00000068; 
    validation_data[  269] = 'h000003aa; 
    validation_data[  270] = 'h000006cf; 
    validation_data[  271] = 'h00000029; 
    validation_data[  272] = 'h000004c3; 
    validation_data[  273] = 'h0000057d; 
    validation_data[  274] = 'h00000791; 
    validation_data[  275] = 'h0000076c; 
    validation_data[  276] = 'h000005fe; 
    validation_data[  277] = 'h00000273; 
    validation_data[  278] = 'h00000153; 
    validation_data[  279] = 'h000004f4; 
    validation_data[  280] = 'h00000691; 
    validation_data[  281] = 'h000003fc; 
    validation_data[  282] = 'h0000028b; 
    validation_data[  283] = 'h0000008f; 
    validation_data[  284] = 'h000006d9; 
    validation_data[  285] = 'h00000024; 
    validation_data[  286] = 'h0000034c; 
    validation_data[  287] = 'h00000628; 
    validation_data[  288] = 'h000003d5; 
    validation_data[  289] = 'h0000065d; 
    validation_data[  290] = 'h000006fa; 
    validation_data[  291] = 'h000006a9; 
    validation_data[  292] = 'h00000170; 
    validation_data[  293] = 'h00000094; 
    validation_data[  294] = 'h00000431; 
    validation_data[  295] = 'h000007ca; 
    validation_data[  296] = 'h00000438; 
    validation_data[  297] = 'h0000063d; 
    validation_data[  298] = 'h0000071b; 
    validation_data[  299] = 'h00000184; 
    validation_data[  300] = 'h000005a5; 
    validation_data[  301] = 'h00000096; 
    validation_data[  302] = 'h0000026f; 
    validation_data[  303] = 'h00000591; 
    validation_data[  304] = 'h0000004e; 
    validation_data[  305] = 'h00000034; 
    validation_data[  306] = 'h0000020c; 
    validation_data[  307] = 'h000001dc; 
    validation_data[  308] = 'h000000bb; 
    validation_data[  309] = 'h0000079f; 
    validation_data[  310] = 'h0000064e; 
    validation_data[  311] = 'h00000693; 
    validation_data[  312] = 'h00000484; 
    validation_data[  313] = 'h00000618; 
    validation_data[  314] = 'h00000776; 
    validation_data[  315] = 'h00000403; 
    validation_data[  316] = 'h000005f6; 
    validation_data[  317] = 'h00000302; 
    validation_data[  318] = 'h000005b1; 
    validation_data[  319] = 'h000004a9; 
    validation_data[  320] = 'h000007e9; 
    validation_data[  321] = 'h000000b8; 
    validation_data[  322] = 'h000006a6; 
    validation_data[  323] = 'h00000726; 
    validation_data[  324] = 'h000002a8; 
    validation_data[  325] = 'h00000438; 
    validation_data[  326] = 'h000001d1; 
    validation_data[  327] = 'h000006fa; 
    validation_data[  328] = 'h0000035b; 
    validation_data[  329] = 'h000000de; 
    validation_data[  330] = 'h000000e4; 
    validation_data[  331] = 'h00000617; 
    validation_data[  332] = 'h000003b1; 
    validation_data[  333] = 'h00000166; 
    validation_data[  334] = 'h00000498; 
    validation_data[  335] = 'h000007e0; 
    validation_data[  336] = 'h0000020c; 
    validation_data[  337] = 'h00000542; 
    validation_data[  338] = 'h00000106; 
    validation_data[  339] = 'h00000559; 
    validation_data[  340] = 'h000003cb; 
    validation_data[  341] = 'h00000366; 
    validation_data[  342] = 'h0000017b; 
    validation_data[  343] = 'h00000750; 
    validation_data[  344] = 'h00000735; 
    validation_data[  345] = 'h000003f2; 
    validation_data[  346] = 'h0000017b; 
    validation_data[  347] = 'h000007e9; 
    validation_data[  348] = 'h000001d3; 
    validation_data[  349] = 'h0000054e; 
    validation_data[  350] = 'h00000098; 
    validation_data[  351] = 'h00000081; 
    validation_data[  352] = 'h00000103; 
    validation_data[  353] = 'h00000547; 
    validation_data[  354] = 'h000006b7; 
    validation_data[  355] = 'h000001b7; 
    validation_data[  356] = 'h00000542; 
    validation_data[  357] = 'h00000729; 
    validation_data[  358] = 'h0000055e; 
    validation_data[  359] = 'h000002ea; 
    validation_data[  360] = 'h00000527; 
    validation_data[  361] = 'h000007d2; 
    validation_data[  362] = 'h000004ed; 
    validation_data[  363] = 'h00000225; 
    validation_data[  364] = 'h000002e9; 
    validation_data[  365] = 'h00000266; 
    validation_data[  366] = 'h00000339; 
    validation_data[  367] = 'h00000277; 
    validation_data[  368] = 'h00000163; 
    validation_data[  369] = 'h0000071d; 
    validation_data[  370] = 'h000007b9; 
    validation_data[  371] = 'h000006a6; 
    validation_data[  372] = 'h00000705; 
    validation_data[  373] = 'h00000553; 
    validation_data[  374] = 'h000000a3; 
    validation_data[  375] = 'h0000062c; 
    validation_data[  376] = 'h00000279; 
    validation_data[  377] = 'h000006f4; 
    validation_data[  378] = 'h00000548; 
    validation_data[  379] = 'h00000313; 
    validation_data[  380] = 'h000005c2; 
    validation_data[  381] = 'h000001b0; 
    validation_data[  382] = 'h000002e7; 
    validation_data[  383] = 'h000000b9; 
    validation_data[  384] = 'h0000033c; 
    validation_data[  385] = 'h000003c7; 
    validation_data[  386] = 'h0000056d; 
    validation_data[  387] = 'h000004bb; 
    validation_data[  388] = 'h00000665; 
    validation_data[  389] = 'h00000115; 
    validation_data[  390] = 'h00000391; 
    validation_data[  391] = 'h0000027b; 
    validation_data[  392] = 'h00000468; 
    validation_data[  393] = 'h000004fc; 
    validation_data[  394] = 'h00000005; 
    validation_data[  395] = 'h000003e1; 
    validation_data[  396] = 'h00000526; 
    validation_data[  397] = 'h000000f1; 
    validation_data[  398] = 'h000002cc; 
    validation_data[  399] = 'h000007e9; 
    validation_data[  400] = 'h0000011f; 
    validation_data[  401] = 'h000004a0; 
    validation_data[  402] = 'h0000072b; 
    validation_data[  403] = 'h0000026f; 
    validation_data[  404] = 'h0000008c; 
    validation_data[  405] = 'h000004ec; 
    validation_data[  406] = 'h00000149; 
    validation_data[  407] = 'h00000248; 
    validation_data[  408] = 'h000001da; 
    validation_data[  409] = 'h000006f8; 
    validation_data[  410] = 'h000002ae; 
    validation_data[  411] = 'h000003a3; 
    validation_data[  412] = 'h0000025f; 
    validation_data[  413] = 'h00000761; 
    validation_data[  414] = 'h00000000; 
    validation_data[  415] = 'h000005e0; 
    validation_data[  416] = 'h000002f5; 
    validation_data[  417] = 'h000001d8; 
    validation_data[  418] = 'h00000225; 
    validation_data[  419] = 'h0000040c; 
    validation_data[  420] = 'h000007a7; 
    validation_data[  421] = 'h00000521; 
    validation_data[  422] = 'h00000617; 
    validation_data[  423] = 'h00000664; 
    validation_data[  424] = 'h000002d3; 
    validation_data[  425] = 'h0000040a; 
    validation_data[  426] = 'h00000398; 
    validation_data[  427] = 'h00000463; 
    validation_data[  428] = 'h00000240; 
    validation_data[  429] = 'h0000018a; 
    validation_data[  430] = 'h000007ad; 
    validation_data[  431] = 'h0000043d; 
    validation_data[  432] = 'h00000487; 
    validation_data[  433] = 'h0000062e; 
    validation_data[  434] = 'h00000003; 
    validation_data[  435] = 'h00000431; 
    validation_data[  436] = 'h000000c3; 
    validation_data[  437] = 'h00000153; 
    validation_data[  438] = 'h000003e1; 
    validation_data[  439] = 'h000000c1; 
    validation_data[  440] = 'h000002a7; 
    validation_data[  441] = 'h0000010e; 
    validation_data[  442] = 'h000001f5; 
    validation_data[  443] = 'h00000396; 
    validation_data[  444] = 'h00000589; 
    validation_data[  445] = 'h00000605; 
    validation_data[  446] = 'h00000307; 
    validation_data[  447] = 'h00000123; 
    validation_data[  448] = 'h00000581; 
    validation_data[  449] = 'h00000527; 
    validation_data[  450] = 'h0000050b; 
    validation_data[  451] = 'h0000038e; 
    validation_data[  452] = 'h00000092; 
    validation_data[  453] = 'h000002ac; 
    validation_data[  454] = 'h000002e1; 
    validation_data[  455] = 'h0000053b; 
    validation_data[  456] = 'h0000062c; 
    validation_data[  457] = 'h000000b6; 
    validation_data[  458] = 'h0000054e; 
    validation_data[  459] = 'h0000027a; 
    validation_data[  460] = 'h000000d7; 
    validation_data[  461] = 'h00000669; 
    validation_data[  462] = 'h0000052e; 
    validation_data[  463] = 'h000002eb; 
    validation_data[  464] = 'h000004db; 
    validation_data[  465] = 'h00000526; 
    validation_data[  466] = 'h00000704; 
    validation_data[  467] = 'h00000508; 
    validation_data[  468] = 'h000004d5; 
    validation_data[  469] = 'h00000690; 
    validation_data[  470] = 'h00000387; 
    validation_data[  471] = 'h00000556; 
    validation_data[  472] = 'h00000398; 
    validation_data[  473] = 'h0000049b; 
    validation_data[  474] = 'h00000640; 
    validation_data[  475] = 'h000004a2; 
    validation_data[  476] = 'h0000003d; 
    validation_data[  477] = 'h000005fd; 
    validation_data[  478] = 'h00000525; 
    validation_data[  479] = 'h000003aa; 
    validation_data[  480] = 'h00000348; 
    validation_data[  481] = 'h000001c8; 
    validation_data[  482] = 'h000000d1; 
    validation_data[  483] = 'h00000479; 
    validation_data[  484] = 'h000002f5; 
    validation_data[  485] = 'h0000044f; 
    validation_data[  486] = 'h000003a3; 
    validation_data[  487] = 'h0000039c; 
    validation_data[  488] = 'h00000175; 
    validation_data[  489] = 'h000001e7; 
    validation_data[  490] = 'h000003e1; 
    validation_data[  491] = 'h000001fc; 
    validation_data[  492] = 'h000003b0; 
    validation_data[  493] = 'h000005ad; 
    validation_data[  494] = 'h00000362; 
    validation_data[  495] = 'h0000061e; 
    validation_data[  496] = 'h00000690; 
    validation_data[  497] = 'h000000da; 
    validation_data[  498] = 'h0000079e; 
    validation_data[  499] = 'h000007fd; 
    validation_data[  500] = 'h000000ea; 
    validation_data[  501] = 'h000006ea; 
    validation_data[  502] = 'h0000028f; 
    validation_data[  503] = 'h00000379; 
    validation_data[  504] = 'h0000073a; 
    validation_data[  505] = 'h00000666; 
    validation_data[  506] = 'h00000500; 
    validation_data[  507] = 'h00000628; 
    validation_data[  508] = 'h00000035; 
    validation_data[  509] = 'h000007d6; 
    validation_data[  510] = 'h000007e2; 
    validation_data[  511] = 'h00000694; 

end


reg clk = 1'b1, rst = 1'b1;
initial #4 rst = 1'b0;
always  #1 clk = ~clk;

wire  miss;
wire [31:0] rd_data;
reg  [31:0] index = 0, wr_data = 0, addr = 0;
reg  rd_req = 1'b0, wr_req = 1'b0;
reg rd_req_ff = 1'b0, miss_ff = 1'b0;
reg [31:0] validation_count = 0;

always @ (posedge clk or posedge rst)
    if(rst) begin
        rd_req_ff <= 1'b0;
        miss_ff   <= 1'b0;
    end else begin
        rd_req_ff <= rd_req;
        miss_ff   <= miss;
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        validation_count <= 0;
    end else begin
        if(validation_count>=`DATA_COUNT) begin
            validation_count <= 'hffffffff;
        end else if(rd_req_ff && (index>(4*`DATA_COUNT))) begin
            if(~miss_ff) begin
                if(validation_data[validation_count]==rd_data)
                    validation_count <= validation_count+1;
                else
                    validation_count <= 0;
            end
        end else begin
            validation_count <= 0;
        end
    end

always @ (posedge clk or posedge rst)
    if(rst) begin
        index   <= 0;
        wr_data <= 0;
        addr    <= 0;
        rd_req  <= 1'b0;
        wr_req  <= 1'b0;
    end else begin
        if(~miss) begin
            if(index<`RDWR_COUNT) begin
                if(wr_cycle[index]) begin
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b1;
                end else if(rd_cycle[index]) begin
                    wr_data <= 0;
                    rd_req  <= 1'b1;
                    wr_req  <= 1'b0;
                end else begin
                    wr_data <= 0;
                    rd_req  <= 1'b0;
                    wr_req  <= 1'b0;
                end
                wr_data <= wr_data_rom[index];
                addr    <= addr_rom[index];
                index <= index + 1;
            end else begin
                wr_data <= 0;
                addr    <= 0;
                rd_req  <= 1'b0;
                wr_req  <= 1'b0;
            end
        end
    end

cache #(
    .LINE_ADDR_LEN  ( 3             ),
    .SET_ADDR_LEN   ( 2             ),
    .TAG_ADDR_LEN   ( 12            ),
    .WAY_CNT        ( 3             )
) cache_test_instance (
    .clk            ( clk           ),
    .rst            ( rst           ),
    .miss           ( miss          ),
    .addr           ( addr          ),
    .rd_req         ( rd_req        ),
    .rd_data        ( rd_data       ),
    .wr_req         ( wr_req        ),
    .wr_data        ( wr_data       )
);

endmodule

