�� 
 m o d u l e   m e m   # (                                       / /    
         p a r a m e t e r     A D D R _ L E N     =   1 1       / /    
 )   (  
         i n p u t     c l k ,   r s t ,  
         i n p u t     [ A D D R _ L E N - 1 : 0 ]   a d d r ,   / /   m e m o r y   a d d r e s s  
         o u t p u t   r e g   [ 3 1 : 0 ]   r d _ d a t a ,     / /   d a t a   r e a d   o u t  
         i n p u t     w r _ r e q ,  
         i n p u t     [ 3 1 : 0 ]   w r _ d a t a               / /   d a t a   w r i t e   i n  
 ) ;  
 l o c a l p a r a m   M E M _ S I Z E   =   1 < < A D D R _ L E N ;  
 r e g   [ 3 1 : 0 ]   r a m _ c e l l   [ M E M _ S I Z E ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )  
                 r d _ d a t a   < =   0 ;  
         e l s e  
                 r d _ d a t a   < =   r a m _ c e l l [ a d d r ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k )  
         i f ( w r _ r e q )    
                 r a m _ c e l l [ a d d r ]   < =   w r _ d a t a ;  
  
 i n i t i a l   b e g i n  
         / /   d s t   m a t r i x   C  
         r a m _ c e l l [               0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 a 1 2 0 8 7 b ;  
         r a m _ c e l l [               1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c a 9 d 7 5 6 b ;  
         r a m _ c e l l [               2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 f e a 4 4 4 f ;  
         r a m _ c e l l [               3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 7 e 2 f 1 0 7 ;  
         r a m _ c e l l [               4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 4 1 a f 7 e 6 ;  
         r a m _ c e l l [               5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 3 f d f 1 c 0 ;  
         r a m _ c e l l [               6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a d c a f d 6 0 ;  
         r a m _ c e l l [               7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 6 0 4 b 6 2 0 ;  
         r a m _ c e l l [               8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 d 5 d 4 f 4 ;  
         r a m _ c e l l [               9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 1 a 9 f 3 7 b ;  
         r a m _ c e l l [             1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 8 8 c d f e 1 ;  
         r a m _ c e l l [             1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 d 2 7 4 d 3 ;  
         r a m _ c e l l [             1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 3 d 9 b f 3 c ;  
         r a m _ c e l l [             1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 1 1 5 6 7 6 c ;  
         r a m _ c e l l [             1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 e 5 1 8 5 8 f ;  
         r a m _ c e l l [             1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 9 0 0 9 f 0 b ;  
         r a m _ c e l l [             1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 0 f 7 2 6 a 0 ;  
         r a m _ c e l l [             1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 a c d b 2 c a ;  
         r a m _ c e l l [             1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 5 d e e 8 1 d ;  
         r a m _ c e l l [             1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a d 3 8 9 6 b 5 ;  
         r a m _ c e l l [             2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 d 2 8 3 0 6 1 ;  
         r a m _ c e l l [             2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 7 7 0 1 5 1 4 ;  
         r a m _ c e l l [             2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 2 4 1 6 5 c 2 ;  
         r a m _ c e l l [             2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 2 b 8 6 c e ;  
         r a m _ c e l l [             2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 b 9 4 7 f 5 5 ;  
         r a m _ c e l l [             2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d e 0 0 1 f 8 5 ;  
         r a m _ c e l l [             2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 7 c c 4 1 e b ;  
         r a m _ c e l l [             2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 b 9 1 1 6 f 9 ;  
         r a m _ c e l l [             2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 0 8 6 b a 5 8 ;  
         r a m _ c e l l [             2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 f 2 6 d 9 8 d ;  
         r a m _ c e l l [             3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 c 2 a f d a 8 ;  
         r a m _ c e l l [             3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 2 a 8 f 9 e ;  
         r a m _ c e l l [             3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e d 7 d b 3 0 c ;  
         r a m _ c e l l [             3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 4 0 5 6 6 9 a ;  
         r a m _ c e l l [             3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 e c f 3 6 b 8 ;  
         r a m _ c e l l [             3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 1 9 8 4 c a 9 ;  
         r a m _ c e l l [             3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e b 3 6 5 9 d f ;  
         r a m _ c e l l [             3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 e 7 1 5 b a b ;  
         r a m _ c e l l [             3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 a c 8 7 2 1 0 ;  
         r a m _ c e l l [             3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b a 6 7 5 9 5 6 ;  
         r a m _ c e l l [             4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 2 6 c 9 a 2 5 ;  
         r a m _ c e l l [             4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 f 0 0 2 2 f b ;  
         r a m _ c e l l [             4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e b 5 2 2 1 3 c ;  
         r a m _ c e l l [             4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 0 9 3 d d 3 ;  
         r a m _ c e l l [             4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b e 2 9 e f e 5 ;  
         r a m _ c e l l [             4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 7 d 5 1 1 e f ;  
         r a m _ c e l l [             4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 4 c 4 8 2 5 9 ;  
         r a m _ c e l l [             4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 6 2 c 4 4 e 4 ;  
         r a m _ c e l l [             4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 b 6 3 c 1 3 d ;  
         r a m _ c e l l [             4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 6 f f 7 a 4 4 ;  
         r a m _ c e l l [             5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f c 6 0 e 7 b d ;  
         r a m _ c e l l [             5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 0 f 9 0 6 6 9 ;  
         r a m _ c e l l [             5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 0 d 4 7 d 2 5 ;  
         r a m _ c e l l [             5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 7 a 8 b e 8 6 ;  
         r a m _ c e l l [             5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 1 9 3 0 8 3 1 ;  
         r a m _ c e l l [             5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 6 b d a 4 a 7 ;  
         r a m _ c e l l [             5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 b 9 6 7 d e f ;  
         r a m _ c e l l [             5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 c f 0 6 3 4 9 ;  
         r a m _ c e l l [             5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 b 8 a e 9 e 5 ;  
         r a m _ c e l l [             5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f a 1 0 7 4 d 3 ;  
         r a m _ c e l l [             6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 5 8 f f e 8 0 ;  
         r a m _ c e l l [             6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 6 e 8 b 6 a 0 ;  
         r a m _ c e l l [             6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 6 1 7 4 b 9 b ;  
         r a m _ c e l l [             6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 6 d 7 4 8 7 8 ;  
         / /   s r c   m a t r i x   A  
         r a m _ c e l l [             6 4 ]   =   3 2 ' h f 9 a 0 d e 8 4 ;  
         r a m _ c e l l [             6 5 ]   =   3 2 ' h d 4 7 7 6 4 d d ;  
         r a m _ c e l l [             6 6 ]   =   3 2 ' h f 4 6 5 a 4 3 7 ;  
         r a m _ c e l l [             6 7 ]   =   3 2 ' h c f 6 6 3 d 7 4 ;  
         r a m _ c e l l [             6 8 ]   =   3 2 ' h f 0 5 d 8 9 e 7 ;  
         r a m _ c e l l [             6 9 ]   =   3 2 ' h a 2 4 3 a 0 4 1 ;  
         r a m _ c e l l [             7 0 ]   =   3 2 ' h a 4 6 5 6 b f 3 ;  
         r a m _ c e l l [             7 1 ]   =   3 2 ' h 8 8 5 0 9 0 e 4 ;  
         r a m _ c e l l [             7 2 ]   =   3 2 ' h 1 0 c a c a f c ;  
         r a m _ c e l l [             7 3 ]   =   3 2 ' h 9 e 3 d 9 f b 8 ;  
         r a m _ c e l l [             7 4 ]   =   3 2 ' h b a 5 2 0 3 3 5 ;  
         r a m _ c e l l [             7 5 ]   =   3 2 ' h b 8 b c 1 3 c d ;  
         r a m _ c e l l [             7 6 ]   =   3 2 ' h 7 2 6 2 9 b e 2 ;  
         r a m _ c e l l [             7 7 ]   =   3 2 ' h b 9 c 2 4 5 8 8 ;  
         r a m _ c e l l [             7 8 ]   =   3 2 ' h 1 b 0 5 7 3 1 3 ;  
         r a m _ c e l l [             7 9 ]   =   3 2 ' h c 9 4 0 a a 9 1 ;  
         r a m _ c e l l [             8 0 ]   =   3 2 ' h 7 9 d 1 f f 5 0 ;  
         r a m _ c e l l [             8 1 ]   =   3 2 ' h 4 f 0 2 b c e a ;  
         r a m _ c e l l [             8 2 ]   =   3 2 ' h 3 d 0 6 f 5 b 1 ;  
         r a m _ c e l l [             8 3 ]   =   3 2 ' h 0 7 4 4 7 6 1 8 ;  
         r a m _ c e l l [             8 4 ]   =   3 2 ' h 9 0 9 b 5 d 5 e ;  
         r a m _ c e l l [             8 5 ]   =   3 2 ' h 6 3 c 6 8 4 a 8 ;  
         r a m _ c e l l [             8 6 ]   =   3 2 ' h 1 5 0 2 d 2 8 3 ;  
         r a m _ c e l l [             8 7 ]   =   3 2 ' h 0 f 2 9 1 f c 1 ;  
         r a m _ c e l l [             8 8 ]   =   3 2 ' h 6 7 1 5 2 b 5 f ;  
         r a m _ c e l l [             8 9 ]   =   3 2 ' h 4 2 b 9 3 7 8 4 ;  
         r a m _ c e l l [             9 0 ]   =   3 2 ' h e b 4 8 c d 5 1 ;  
         r a m _ c e l l [             9 1 ]   =   3 2 ' h f 7 b 7 0 e 6 b ;  
         r a m _ c e l l [             9 2 ]   =   3 2 ' h f 9 f b 9 7 d 5 ;  
         r a m _ c e l l [             9 3 ]   =   3 2 ' h d 3 5 0 1 f 6 8 ;  
         r a m _ c e l l [             9 4 ]   =   3 2 ' h 6 b f 8 4 7 a 6 ;  
         r a m _ c e l l [             9 5 ]   =   3 2 ' h c e 9 c 4 a 9 c ;  
         r a m _ c e l l [             9 6 ]   =   3 2 ' h e e 3 9 7 e f 3 ;  
         r a m _ c e l l [             9 7 ]   =   3 2 ' h 2 5 3 7 7 9 5 9 ;  
         r a m _ c e l l [             9 8 ]   =   3 2 ' h 1 9 f 1 4 4 d e ;  
         r a m _ c e l l [             9 9 ]   =   3 2 ' h 3 5 f 6 0 7 d 6 ;  
         r a m _ c e l l [           1 0 0 ]   =   3 2 ' h 8 5 8 8 9 1 9 e ;  
         r a m _ c e l l [           1 0 1 ]   =   3 2 ' h 4 a 9 4 a 7 d e ;  
         r a m _ c e l l [           1 0 2 ]   =   3 2 ' h 7 d 5 d b 4 4 b ;  
         r a m _ c e l l [           1 0 3 ]   =   3 2 ' h 1 b 8 7 b 7 a a ;  
         r a m _ c e l l [           1 0 4 ]   =   3 2 ' h 9 4 b a b 5 7 7 ;  
         r a m _ c e l l [           1 0 5 ]   =   3 2 ' h 5 5 7 0 e 4 e 6 ;  
         r a m _ c e l l [           1 0 6 ]   =   3 2 ' h d 6 6 e 1 b 3 e ;  
         r a m _ c e l l [           1 0 7 ]   =   3 2 ' h 6 8 5 9 8 f 0 7 ;  
         r a m _ c e l l [           1 0 8 ]   =   3 2 ' h 6 3 b b a 4 e 3 ;  
         r a m _ c e l l [           1 0 9 ]   =   3 2 ' h d b 2 0 a d 4 b ;  
         r a m _ c e l l [           1 1 0 ]   =   3 2 ' h 7 d 0 5 7 e 2 5 ;  
         r a m _ c e l l [           1 1 1 ]   =   3 2 ' h f 1 3 9 9 b 7 8 ;  
         r a m _ c e l l [           1 1 2 ]   =   3 2 ' h e b 6 7 e b c d ;  
         r a m _ c e l l [           1 1 3 ]   =   3 2 ' h e 8 2 5 3 4 3 f ;  
         r a m _ c e l l [           1 1 4 ]   =   3 2 ' h 9 7 7 f 7 a d 0 ;  
         r a m _ c e l l [           1 1 5 ]   =   3 2 ' h 9 6 8 4 1 b 4 0 ;  
         r a m _ c e l l [           1 1 6 ]   =   3 2 ' h 6 d 2 c d c 2 b ;  
         r a m _ c e l l [           1 1 7 ]   =   3 2 ' h c b 2 3 d 6 0 9 ;  
         r a m _ c e l l [           1 1 8 ]   =   3 2 ' h 8 c 4 4 8 8 d 1 ;  
         r a m _ c e l l [           1 1 9 ]   =   3 2 ' h 1 e 6 c 0 6 c 5 ;  
         r a m _ c e l l [           1 2 0 ]   =   3 2 ' h 0 7 c 8 8 a a 2 ;  
         r a m _ c e l l [           1 2 1 ]   =   3 2 ' h c 8 5 a e c e a ;  
         r a m _ c e l l [           1 2 2 ]   =   3 2 ' h c c d 1 b d 6 1 ;  
         r a m _ c e l l [           1 2 3 ]   =   3 2 ' h f 9 f 1 5 a c c ;  
         r a m _ c e l l [           1 2 4 ]   =   3 2 ' h 7 e e 3 4 7 3 d ;  
         r a m _ c e l l [           1 2 5 ]   =   3 2 ' h 5 7 e 7 9 e 7 6 ;  
         r a m _ c e l l [           1 2 6 ]   =   3 2 ' h e f e 7 5 2 e a ;  
         r a m _ c e l l [           1 2 7 ]   =   3 2 ' h 4 1 2 2 b 2 7 3 ;  
         / /   s r c   m a t r i x   B  
         r a m _ c e l l [           1 2 8 ]   =   3 2 ' h a a 1 e d 8 e 8 ;  
         r a m _ c e l l [           1 2 9 ]   =   3 2 ' h b 2 b e 3 1 2 0 ;  
         r a m _ c e l l [           1 3 0 ]   =   3 2 ' h 5 9 1 7 0 f 5 c ;  
         r a m _ c e l l [           1 3 1 ]   =   3 2 ' h f d d 6 d 2 2 4 ;  
         r a m _ c e l l [           1 3 2 ]   =   3 2 ' h 9 f b 3 1 5 9 d ;  
         r a m _ c e l l [           1 3 3 ]   =   3 2 ' h 0 d c 2 d 2 8 1 ;  
         r a m _ c e l l [           1 3 4 ]   =   3 2 ' h 0 c 3 9 f b 3 2 ;  
         r a m _ c e l l [           1 3 5 ]   =   3 2 ' h e 4 b a 4 7 7 e ;  
         r a m _ c e l l [           1 3 6 ]   =   3 2 ' h 6 a d 3 c 5 d 4 ;  
         r a m _ c e l l [           1 3 7 ]   =   3 2 ' h 2 1 6 a 9 2 5 5 ;  
         r a m _ c e l l [           1 3 8 ]   =   3 2 ' h e 9 1 d c a c 5 ;  
         r a m _ c e l l [           1 3 9 ]   =   3 2 ' h 7 a d 6 5 e 3 a ;  
         r a m _ c e l l [           1 4 0 ]   =   3 2 ' h 9 3 e 6 c 2 d 7 ;  
         r a m _ c e l l [           1 4 1 ]   =   3 2 ' h 3 f d 4 7 b 4 d ;  
         r a m _ c e l l [           1 4 2 ]   =   3 2 ' h 8 3 1 6 3 9 7 1 ;  
         r a m _ c e l l [           1 4 3 ]   =   3 2 ' h 8 6 c 4 d b 7 9 ;  
         r a m _ c e l l [           1 4 4 ]   =   3 2 ' h 0 1 a f d f 3 6 ;  
         r a m _ c e l l [           1 4 5 ]   =   3 2 ' h 3 f 5 f d 1 a 8 ;  
         r a m _ c e l l [           1 4 6 ]   =   3 2 ' h 0 f 5 e 0 5 3 8 ;  
         r a m _ c e l l [           1 4 7 ]   =   3 2 ' h 2 c 3 5 f 8 d 6 ;  
         r a m _ c e l l [           1 4 8 ]   =   3 2 ' h 2 b f e c 8 d e ;  
         r a m _ c e l l [           1 4 9 ]   =   3 2 ' h 6 e c 5 6 3 7 7 ;  
         r a m _ c e l l [           1 5 0 ]   =   3 2 ' h c 8 b 7 d 2 6 9 ;  
         r a m _ c e l l [           1 5 1 ]   =   3 2 ' h d 4 c 0 2 0 3 4 ;  
         r a m _ c e l l [           1 5 2 ]   =   3 2 ' h d d 1 3 8 d 7 0 ;  
         r a m _ c e l l [           1 5 3 ]   =   3 2 ' h f 2 e 2 d 9 5 1 ;  
         r a m _ c e l l [           1 5 4 ]   =   3 2 ' h 8 3 7 5 e 6 a 0 ;  
         r a m _ c e l l [           1 5 5 ]   =   3 2 ' h 3 3 4 5 5 a 2 2 ;  
         r a m _ c e l l [           1 5 6 ]   =   3 2 ' h d 9 9 9 3 8 0 9 ;  
         r a m _ c e l l [           1 5 7 ]   =   3 2 ' h 8 f b f 9 b d e ;  
         r a m _ c e l l [           1 5 8 ]   =   3 2 ' h 5 9 2 3 0 0 9 3 ;  
         r a m _ c e l l [           1 5 9 ]   =   3 2 ' h 4 6 8 8 e 6 8 d ;  
         r a m _ c e l l [           1 6 0 ]   =   3 2 ' h b f f 3 2 2 9 9 ;  
         r a m _ c e l l [           1 6 1 ]   =   3 2 ' h e 3 0 d 4 6 f 0 ;  
         r a m _ c e l l [           1 6 2 ]   =   3 2 ' h 2 a 7 5 5 b d b ;  
         r a m _ c e l l [           1 6 3 ]   =   3 2 ' h c 1 f f 4 3 5 9 ;  
         r a m _ c e l l [           1 6 4 ]   =   3 2 ' h b 7 8 b d 2 7 4 ;  
         r a m _ c e l l [           1 6 5 ]   =   3 2 ' h 9 a 9 f 4 7 e 3 ;  
         r a m _ c e l l [           1 6 6 ]   =   3 2 ' h 9 d 1 9 8 1 f 6 ;  
         r a m _ c e l l [           1 6 7 ]   =   3 2 ' h 5 5 e a 5 6 9 b ;  
         r a m _ c e l l [           1 6 8 ]   =   3 2 ' h 0 1 4 8 0 7 9 e ;  
         r a m _ c e l l [           1 6 9 ]   =   3 2 ' h 3 7 f 1 b 0 d 9 ;  
         r a m _ c e l l [           1 7 0 ]   =   3 2 ' h a b 6 e a a 8 0 ;  
         r a m _ c e l l [           1 7 1 ]   =   3 2 ' h 2 6 9 8 7 e b 7 ;  
         r a m _ c e l l [           1 7 2 ]   =   3 2 ' h 5 8 1 2 6 a 7 6 ;  
         r a m _ c e l l [           1 7 3 ]   =   3 2 ' h f b 0 8 2 6 0 2 ;  
         r a m _ c e l l [           1 7 4 ]   =   3 2 ' h 9 c 3 5 3 7 d 9 ;  
         r a m _ c e l l [           1 7 5 ]   =   3 2 ' h 4 2 3 e d 0 1 5 ;  
         r a m _ c e l l [           1 7 6 ]   =   3 2 ' h f 7 9 d d c c 0 ;  
         r a m _ c e l l [           1 7 7 ]   =   3 2 ' h a 2 f f 2 9 e d ;  
         r a m _ c e l l [           1 7 8 ]   =   3 2 ' h 8 5 d f 2 3 5 b ;  
         r a m _ c e l l [           1 7 9 ]   =   3 2 ' h 3 6 5 d 1 0 d b ;  
         r a m _ c e l l [           1 8 0 ]   =   3 2 ' h f 3 e 4 5 9 3 b ;  
         r a m _ c e l l [           1 8 1 ]   =   3 2 ' h 6 3 f a 6 3 2 9 ;  
         r a m _ c e l l [           1 8 2 ]   =   3 2 ' h d f 2 1 7 0 7 3 ;  
         r a m _ c e l l [           1 8 3 ]   =   3 2 ' h 7 4 c d 6 a c 3 ;  
         r a m _ c e l l [           1 8 4 ]   =   3 2 ' h 1 2 0 9 7 b 4 0 ;  
         r a m _ c e l l [           1 8 5 ]   =   3 2 ' h 8 6 e a 2 a a 5 ;  
         r a m _ c e l l [           1 8 6 ]   =   3 2 ' h e b f b 0 9 2 a ;  
         r a m _ c e l l [           1 8 7 ]   =   3 2 ' h a 3 8 7 2 f b 0 ;  
         r a m _ c e l l [           1 8 8 ]   =   3 2 ' h e 5 c 2 0 9 a a ;  
         r a m _ c e l l [           1 8 9 ]   =   3 2 ' h 7 7 4 d 0 c 6 c ;  
         r a m _ c e l l [           1 9 0 ]   =   3 2 ' h a 9 9 f a c 5 6 ;  
         r a m _ c e l l [           1 9 1 ]   =   3 2 ' h 0 1 5 9 0 a 5 7 ;  
 e n d  
  
 e n d m o d u l e  
  
 