
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h4b81cb67;
    ram_cell[       1] = 32'h0;  // 32'haa597913;
    ram_cell[       2] = 32'h0;  // 32'h5eb89271;
    ram_cell[       3] = 32'h0;  // 32'h4173350f;
    ram_cell[       4] = 32'h0;  // 32'h4c21436f;
    ram_cell[       5] = 32'h0;  // 32'h41bc852c;
    ram_cell[       6] = 32'h0;  // 32'h603eba11;
    ram_cell[       7] = 32'h0;  // 32'h63801ec3;
    ram_cell[       8] = 32'h0;  // 32'ha86b321e;
    ram_cell[       9] = 32'h0;  // 32'h70748bd0;
    ram_cell[      10] = 32'h0;  // 32'h438140ae;
    ram_cell[      11] = 32'h0;  // 32'h2ac82cc3;
    ram_cell[      12] = 32'h0;  // 32'h0f7ed628;
    ram_cell[      13] = 32'h0;  // 32'h3a624755;
    ram_cell[      14] = 32'h0;  // 32'h7282c0f6;
    ram_cell[      15] = 32'h0;  // 32'h78676d2b;
    ram_cell[      16] = 32'h0;  // 32'h18b95249;
    ram_cell[      17] = 32'h0;  // 32'hd75d8e55;
    ram_cell[      18] = 32'h0;  // 32'h454e0585;
    ram_cell[      19] = 32'h0;  // 32'hd22b17f1;
    ram_cell[      20] = 32'h0;  // 32'ha8102849;
    ram_cell[      21] = 32'h0;  // 32'hb1eed3e9;
    ram_cell[      22] = 32'h0;  // 32'h17c6043a;
    ram_cell[      23] = 32'h0;  // 32'h65ef040d;
    ram_cell[      24] = 32'h0;  // 32'ha0bcdb00;
    ram_cell[      25] = 32'h0;  // 32'h85d9e975;
    ram_cell[      26] = 32'h0;  // 32'h362bd763;
    ram_cell[      27] = 32'h0;  // 32'h55922d78;
    ram_cell[      28] = 32'h0;  // 32'hd05872c6;
    ram_cell[      29] = 32'h0;  // 32'heb96fd91;
    ram_cell[      30] = 32'h0;  // 32'h73916ed5;
    ram_cell[      31] = 32'h0;  // 32'h044aa44a;
    ram_cell[      32] = 32'h0;  // 32'hf7ca0057;
    ram_cell[      33] = 32'h0;  // 32'h427b1df9;
    ram_cell[      34] = 32'h0;  // 32'hd1ab0af8;
    ram_cell[      35] = 32'h0;  // 32'hb1808f5b;
    ram_cell[      36] = 32'h0;  // 32'hf6fc94c2;
    ram_cell[      37] = 32'h0;  // 32'h132c8233;
    ram_cell[      38] = 32'h0;  // 32'h51f62a8c;
    ram_cell[      39] = 32'h0;  // 32'hd610dae9;
    ram_cell[      40] = 32'h0;  // 32'h93abbd28;
    ram_cell[      41] = 32'h0;  // 32'hbb3ad2b7;
    ram_cell[      42] = 32'h0;  // 32'h0682b6cb;
    ram_cell[      43] = 32'h0;  // 32'hcb999438;
    ram_cell[      44] = 32'h0;  // 32'hf3c3f426;
    ram_cell[      45] = 32'h0;  // 32'ha336cae3;
    ram_cell[      46] = 32'h0;  // 32'h537ec3cd;
    ram_cell[      47] = 32'h0;  // 32'h3ec5c1ed;
    ram_cell[      48] = 32'h0;  // 32'h5fd2d00f;
    ram_cell[      49] = 32'h0;  // 32'h2239e5ae;
    ram_cell[      50] = 32'h0;  // 32'hda3577f1;
    ram_cell[      51] = 32'h0;  // 32'h69341e31;
    ram_cell[      52] = 32'h0;  // 32'hc448e948;
    ram_cell[      53] = 32'h0;  // 32'h0d9a69ae;
    ram_cell[      54] = 32'h0;  // 32'h3feea8af;
    ram_cell[      55] = 32'h0;  // 32'h01bc1036;
    ram_cell[      56] = 32'h0;  // 32'h1feefbbb;
    ram_cell[      57] = 32'h0;  // 32'h2b9fcbe9;
    ram_cell[      58] = 32'h0;  // 32'hda45f0d0;
    ram_cell[      59] = 32'h0;  // 32'hfd9473aa;
    ram_cell[      60] = 32'h0;  // 32'hfe46ee20;
    ram_cell[      61] = 32'h0;  // 32'hfa4067e6;
    ram_cell[      62] = 32'h0;  // 32'h0f8c4f19;
    ram_cell[      63] = 32'h0;  // 32'he233ed08;
    ram_cell[      64] = 32'h0;  // 32'h861ca3d8;
    ram_cell[      65] = 32'h0;  // 32'ha6753f32;
    ram_cell[      66] = 32'h0;  // 32'h15b329eb;
    ram_cell[      67] = 32'h0;  // 32'h241ce5b6;
    ram_cell[      68] = 32'h0;  // 32'hebc98ea5;
    ram_cell[      69] = 32'h0;  // 32'h9260cb68;
    ram_cell[      70] = 32'h0;  // 32'h15c286c1;
    ram_cell[      71] = 32'h0;  // 32'h3dae70c6;
    ram_cell[      72] = 32'h0;  // 32'hc6a8ee41;
    ram_cell[      73] = 32'h0;  // 32'h8b84da00;
    ram_cell[      74] = 32'h0;  // 32'h9e124804;
    ram_cell[      75] = 32'h0;  // 32'h5fb8c663;
    ram_cell[      76] = 32'h0;  // 32'h6d95d188;
    ram_cell[      77] = 32'h0;  // 32'hce89d648;
    ram_cell[      78] = 32'h0;  // 32'h45e45eea;
    ram_cell[      79] = 32'h0;  // 32'hd794dfa4;
    ram_cell[      80] = 32'h0;  // 32'h407a4dee;
    ram_cell[      81] = 32'h0;  // 32'hfa56267e;
    ram_cell[      82] = 32'h0;  // 32'h19ca0d51;
    ram_cell[      83] = 32'h0;  // 32'h9fefa42f;
    ram_cell[      84] = 32'h0;  // 32'hae4f9859;
    ram_cell[      85] = 32'h0;  // 32'h97e4ded9;
    ram_cell[      86] = 32'h0;  // 32'h32c1e474;
    ram_cell[      87] = 32'h0;  // 32'h0ae5f229;
    ram_cell[      88] = 32'h0;  // 32'h04de74b7;
    ram_cell[      89] = 32'h0;  // 32'h16c2c15d;
    ram_cell[      90] = 32'h0;  // 32'hd27ca753;
    ram_cell[      91] = 32'h0;  // 32'h2aedfa40;
    ram_cell[      92] = 32'h0;  // 32'h8716f0f7;
    ram_cell[      93] = 32'h0;  // 32'hd5d3133b;
    ram_cell[      94] = 32'h0;  // 32'h5c2b4840;
    ram_cell[      95] = 32'h0;  // 32'he0ebe4d0;
    ram_cell[      96] = 32'h0;  // 32'h2dc8be03;
    ram_cell[      97] = 32'h0;  // 32'hb9964578;
    ram_cell[      98] = 32'h0;  // 32'hba4bf668;
    ram_cell[      99] = 32'h0;  // 32'h86bd4e46;
    ram_cell[     100] = 32'h0;  // 32'h7fb91527;
    ram_cell[     101] = 32'h0;  // 32'h2840c796;
    ram_cell[     102] = 32'h0;  // 32'h6052cc98;
    ram_cell[     103] = 32'h0;  // 32'h6b5546b3;
    ram_cell[     104] = 32'h0;  // 32'h772c45ad;
    ram_cell[     105] = 32'h0;  // 32'h9fb6424f;
    ram_cell[     106] = 32'h0;  // 32'h7724694d;
    ram_cell[     107] = 32'h0;  // 32'hd7c61e56;
    ram_cell[     108] = 32'h0;  // 32'h5ce99708;
    ram_cell[     109] = 32'h0;  // 32'h8be1f29b;
    ram_cell[     110] = 32'h0;  // 32'hea7524e9;
    ram_cell[     111] = 32'h0;  // 32'h5aa8b972;
    ram_cell[     112] = 32'h0;  // 32'h5f1fe799;
    ram_cell[     113] = 32'h0;  // 32'h4d945ea3;
    ram_cell[     114] = 32'h0;  // 32'ha571e0ed;
    ram_cell[     115] = 32'h0;  // 32'h9dead70a;
    ram_cell[     116] = 32'h0;  // 32'h05032b0e;
    ram_cell[     117] = 32'h0;  // 32'hc4260795;
    ram_cell[     118] = 32'h0;  // 32'h7b894b2b;
    ram_cell[     119] = 32'h0;  // 32'he7fa84f2;
    ram_cell[     120] = 32'h0;  // 32'hca6b92c1;
    ram_cell[     121] = 32'h0;  // 32'h57d466ad;
    ram_cell[     122] = 32'h0;  // 32'hda60ba54;
    ram_cell[     123] = 32'h0;  // 32'h9893fcdc;
    ram_cell[     124] = 32'h0;  // 32'h30a2e59d;
    ram_cell[     125] = 32'h0;  // 32'h9d65f29a;
    ram_cell[     126] = 32'h0;  // 32'h63222c6c;
    ram_cell[     127] = 32'h0;  // 32'hef9c8ea5;
    ram_cell[     128] = 32'h0;  // 32'ha3ebf081;
    ram_cell[     129] = 32'h0;  // 32'h55c3fb64;
    ram_cell[     130] = 32'h0;  // 32'hc176213a;
    ram_cell[     131] = 32'h0;  // 32'h53355b66;
    ram_cell[     132] = 32'h0;  // 32'ha5059c8a;
    ram_cell[     133] = 32'h0;  // 32'hbc9d8416;
    ram_cell[     134] = 32'h0;  // 32'hf1c4eaae;
    ram_cell[     135] = 32'h0;  // 32'h52b41de0;
    ram_cell[     136] = 32'h0;  // 32'h965560f7;
    ram_cell[     137] = 32'h0;  // 32'h81605271;
    ram_cell[     138] = 32'h0;  // 32'h324c1957;
    ram_cell[     139] = 32'h0;  // 32'hc3ff916a;
    ram_cell[     140] = 32'h0;  // 32'h62ad1ebe;
    ram_cell[     141] = 32'h0;  // 32'h518339a4;
    ram_cell[     142] = 32'h0;  // 32'h37d9f2f2;
    ram_cell[     143] = 32'h0;  // 32'hcfe2825f;
    ram_cell[     144] = 32'h0;  // 32'h0c73f1a8;
    ram_cell[     145] = 32'h0;  // 32'hc9838673;
    ram_cell[     146] = 32'h0;  // 32'hac5e619a;
    ram_cell[     147] = 32'h0;  // 32'hdd244b08;
    ram_cell[     148] = 32'h0;  // 32'h20e5c4ae;
    ram_cell[     149] = 32'h0;  // 32'h975bea1d;
    ram_cell[     150] = 32'h0;  // 32'h387f1fe2;
    ram_cell[     151] = 32'h0;  // 32'hefdb3555;
    ram_cell[     152] = 32'h0;  // 32'h43c89110;
    ram_cell[     153] = 32'h0;  // 32'he6ac2112;
    ram_cell[     154] = 32'h0;  // 32'hd016ae2f;
    ram_cell[     155] = 32'h0;  // 32'h649354bd;
    ram_cell[     156] = 32'h0;  // 32'h632ae8b2;
    ram_cell[     157] = 32'h0;  // 32'haeb28fec;
    ram_cell[     158] = 32'h0;  // 32'h9472123c;
    ram_cell[     159] = 32'h0;  // 32'h60665964;
    ram_cell[     160] = 32'h0;  // 32'h279d8bf0;
    ram_cell[     161] = 32'h0;  // 32'h2131263e;
    ram_cell[     162] = 32'h0;  // 32'h10fdb0ba;
    ram_cell[     163] = 32'h0;  // 32'h4bd030dd;
    ram_cell[     164] = 32'h0;  // 32'hcf84df69;
    ram_cell[     165] = 32'h0;  // 32'hd0d3e942;
    ram_cell[     166] = 32'h0;  // 32'hbeb0d680;
    ram_cell[     167] = 32'h0;  // 32'h71574b77;
    ram_cell[     168] = 32'h0;  // 32'he2494b0c;
    ram_cell[     169] = 32'h0;  // 32'hee2380a4;
    ram_cell[     170] = 32'h0;  // 32'hb36d2b31;
    ram_cell[     171] = 32'h0;  // 32'h1426bafc;
    ram_cell[     172] = 32'h0;  // 32'h6916df19;
    ram_cell[     173] = 32'h0;  // 32'hf90cc268;
    ram_cell[     174] = 32'h0;  // 32'hded8f9e4;
    ram_cell[     175] = 32'h0;  // 32'h684597db;
    ram_cell[     176] = 32'h0;  // 32'h52a24d85;
    ram_cell[     177] = 32'h0;  // 32'hc0c0f4d8;
    ram_cell[     178] = 32'h0;  // 32'h5c478b02;
    ram_cell[     179] = 32'h0;  // 32'h36a21c22;
    ram_cell[     180] = 32'h0;  // 32'h1bc99c3c;
    ram_cell[     181] = 32'h0;  // 32'h213b9ad4;
    ram_cell[     182] = 32'h0;  // 32'h6301d2d1;
    ram_cell[     183] = 32'h0;  // 32'haff88481;
    ram_cell[     184] = 32'h0;  // 32'h855277e5;
    ram_cell[     185] = 32'h0;  // 32'h5336afa7;
    ram_cell[     186] = 32'h0;  // 32'h97e67d39;
    ram_cell[     187] = 32'h0;  // 32'h5995a423;
    ram_cell[     188] = 32'h0;  // 32'hebd49718;
    ram_cell[     189] = 32'h0;  // 32'h6fc37259;
    ram_cell[     190] = 32'h0;  // 32'h4f836e59;
    ram_cell[     191] = 32'h0;  // 32'h5b88b078;
    ram_cell[     192] = 32'h0;  // 32'he92111a8;
    ram_cell[     193] = 32'h0;  // 32'hbc9ce608;
    ram_cell[     194] = 32'h0;  // 32'h34cf13b8;
    ram_cell[     195] = 32'h0;  // 32'h685b1738;
    ram_cell[     196] = 32'h0;  // 32'hb6c3b339;
    ram_cell[     197] = 32'h0;  // 32'h32a4f9f6;
    ram_cell[     198] = 32'h0;  // 32'hcf312c46;
    ram_cell[     199] = 32'h0;  // 32'h5fa893aa;
    ram_cell[     200] = 32'h0;  // 32'h28eea390;
    ram_cell[     201] = 32'h0;  // 32'h5e602636;
    ram_cell[     202] = 32'h0;  // 32'hc6d6b3a5;
    ram_cell[     203] = 32'h0;  // 32'h3912cd8c;
    ram_cell[     204] = 32'h0;  // 32'h47754287;
    ram_cell[     205] = 32'h0;  // 32'hbbe0a2f2;
    ram_cell[     206] = 32'h0;  // 32'h4b57598a;
    ram_cell[     207] = 32'h0;  // 32'h0235ed75;
    ram_cell[     208] = 32'h0;  // 32'he08a8ac6;
    ram_cell[     209] = 32'h0;  // 32'h512d031b;
    ram_cell[     210] = 32'h0;  // 32'h2a98906c;
    ram_cell[     211] = 32'h0;  // 32'h308c3b91;
    ram_cell[     212] = 32'h0;  // 32'h778d7712;
    ram_cell[     213] = 32'h0;  // 32'hfb6cb553;
    ram_cell[     214] = 32'h0;  // 32'h2f1382e3;
    ram_cell[     215] = 32'h0;  // 32'h2e666414;
    ram_cell[     216] = 32'h0;  // 32'h4d6f3e1c;
    ram_cell[     217] = 32'h0;  // 32'h6e0cb16c;
    ram_cell[     218] = 32'h0;  // 32'h43fe28ed;
    ram_cell[     219] = 32'h0;  // 32'h6252e126;
    ram_cell[     220] = 32'h0;  // 32'h9e60a706;
    ram_cell[     221] = 32'h0;  // 32'he47ce87e;
    ram_cell[     222] = 32'h0;  // 32'hd2d54790;
    ram_cell[     223] = 32'h0;  // 32'h2ae8366d;
    ram_cell[     224] = 32'h0;  // 32'h372b4274;
    ram_cell[     225] = 32'h0;  // 32'h7c665e3d;
    ram_cell[     226] = 32'h0;  // 32'h4e2c79bb;
    ram_cell[     227] = 32'h0;  // 32'h3a3d14b5;
    ram_cell[     228] = 32'h0;  // 32'hd88af11f;
    ram_cell[     229] = 32'h0;  // 32'h50fe43e9;
    ram_cell[     230] = 32'h0;  // 32'h50851ebf;
    ram_cell[     231] = 32'h0;  // 32'hf447d165;
    ram_cell[     232] = 32'h0;  // 32'h28f8acaa;
    ram_cell[     233] = 32'h0;  // 32'h4e6b945e;
    ram_cell[     234] = 32'h0;  // 32'hafcf6a9a;
    ram_cell[     235] = 32'h0;  // 32'h0c153dda;
    ram_cell[     236] = 32'h0;  // 32'h17f3e3cf;
    ram_cell[     237] = 32'h0;  // 32'h49874850;
    ram_cell[     238] = 32'h0;  // 32'hb49d1229;
    ram_cell[     239] = 32'h0;  // 32'h3f21a240;
    ram_cell[     240] = 32'h0;  // 32'hd91c4ad9;
    ram_cell[     241] = 32'h0;  // 32'h6b0a38b8;
    ram_cell[     242] = 32'h0;  // 32'h2a7cf7bd;
    ram_cell[     243] = 32'h0;  // 32'h147e43d9;
    ram_cell[     244] = 32'h0;  // 32'h09e1ea52;
    ram_cell[     245] = 32'h0;  // 32'h62df2b57;
    ram_cell[     246] = 32'h0;  // 32'hf60118bc;
    ram_cell[     247] = 32'h0;  // 32'had1bce2f;
    ram_cell[     248] = 32'h0;  // 32'h7c11ce1e;
    ram_cell[     249] = 32'h0;  // 32'hc5dd8b52;
    ram_cell[     250] = 32'h0;  // 32'h644a2370;
    ram_cell[     251] = 32'h0;  // 32'h14abba65;
    ram_cell[     252] = 32'h0;  // 32'h542c6049;
    ram_cell[     253] = 32'h0;  // 32'hef51d282;
    ram_cell[     254] = 32'h0;  // 32'h49dbe5c3;
    ram_cell[     255] = 32'h0;  // 32'h0eb46165;
    // src matrix A
    ram_cell[     256] = 32'hb6b03bf9;
    ram_cell[     257] = 32'h699ec11f;
    ram_cell[     258] = 32'hf3b8b62f;
    ram_cell[     259] = 32'h89726e1d;
    ram_cell[     260] = 32'h2e3fccae;
    ram_cell[     261] = 32'h3c920811;
    ram_cell[     262] = 32'h8cf23d19;
    ram_cell[     263] = 32'h58b8e710;
    ram_cell[     264] = 32'hbc0854a4;
    ram_cell[     265] = 32'hec99df41;
    ram_cell[     266] = 32'h7ef18f89;
    ram_cell[     267] = 32'hdf7e2383;
    ram_cell[     268] = 32'h5a2a7800;
    ram_cell[     269] = 32'hebf2cfea;
    ram_cell[     270] = 32'hb04b1a67;
    ram_cell[     271] = 32'h365f870b;
    ram_cell[     272] = 32'h8c958fc1;
    ram_cell[     273] = 32'h28e7772f;
    ram_cell[     274] = 32'h445c4674;
    ram_cell[     275] = 32'h9a953f23;
    ram_cell[     276] = 32'h63cd4d07;
    ram_cell[     277] = 32'hf8e6c590;
    ram_cell[     278] = 32'h001de0c1;
    ram_cell[     279] = 32'h015d8111;
    ram_cell[     280] = 32'hc7641fb0;
    ram_cell[     281] = 32'h1f91a4bd;
    ram_cell[     282] = 32'h9cf151bd;
    ram_cell[     283] = 32'h297accad;
    ram_cell[     284] = 32'h30d54114;
    ram_cell[     285] = 32'h3a35295c;
    ram_cell[     286] = 32'h3c264d7e;
    ram_cell[     287] = 32'h77c19c04;
    ram_cell[     288] = 32'hd8144545;
    ram_cell[     289] = 32'h8b28bb58;
    ram_cell[     290] = 32'h7bc94a33;
    ram_cell[     291] = 32'h634f507e;
    ram_cell[     292] = 32'h8b3bf1c7;
    ram_cell[     293] = 32'hb952c155;
    ram_cell[     294] = 32'he9ac4895;
    ram_cell[     295] = 32'h3491a394;
    ram_cell[     296] = 32'h5bc9bd43;
    ram_cell[     297] = 32'ha33d3dd6;
    ram_cell[     298] = 32'had9edf03;
    ram_cell[     299] = 32'h5288f1b9;
    ram_cell[     300] = 32'hda6bc2f0;
    ram_cell[     301] = 32'ha09bded1;
    ram_cell[     302] = 32'he3b326b5;
    ram_cell[     303] = 32'h6fa737c9;
    ram_cell[     304] = 32'h4dcee6a2;
    ram_cell[     305] = 32'hb353b741;
    ram_cell[     306] = 32'h76b0ea66;
    ram_cell[     307] = 32'h5aac90d0;
    ram_cell[     308] = 32'h8180600f;
    ram_cell[     309] = 32'h97d842fb;
    ram_cell[     310] = 32'h08a03371;
    ram_cell[     311] = 32'he01f8ff7;
    ram_cell[     312] = 32'h6197b487;
    ram_cell[     313] = 32'hd2b22011;
    ram_cell[     314] = 32'h6f7b7a47;
    ram_cell[     315] = 32'h18385769;
    ram_cell[     316] = 32'h82abb6df;
    ram_cell[     317] = 32'hca752abc;
    ram_cell[     318] = 32'h4a47de8d;
    ram_cell[     319] = 32'h695b68f6;
    ram_cell[     320] = 32'h104530de;
    ram_cell[     321] = 32'h33c6e9c1;
    ram_cell[     322] = 32'hf3e0116a;
    ram_cell[     323] = 32'h9ee9e567;
    ram_cell[     324] = 32'h3e2681f2;
    ram_cell[     325] = 32'h1bf31b69;
    ram_cell[     326] = 32'h7f19a19a;
    ram_cell[     327] = 32'hf9118089;
    ram_cell[     328] = 32'h9481432c;
    ram_cell[     329] = 32'h1554d458;
    ram_cell[     330] = 32'h8e4f5d9d;
    ram_cell[     331] = 32'h92d6eeef;
    ram_cell[     332] = 32'h921f659a;
    ram_cell[     333] = 32'h109cd919;
    ram_cell[     334] = 32'h32592f23;
    ram_cell[     335] = 32'h5591994d;
    ram_cell[     336] = 32'h46528b89;
    ram_cell[     337] = 32'hdd3acac8;
    ram_cell[     338] = 32'h3e44f674;
    ram_cell[     339] = 32'h056dd752;
    ram_cell[     340] = 32'h9433617f;
    ram_cell[     341] = 32'h6f56a6c5;
    ram_cell[     342] = 32'ha2fca485;
    ram_cell[     343] = 32'hc29d8965;
    ram_cell[     344] = 32'hbc18525c;
    ram_cell[     345] = 32'hd5c7f507;
    ram_cell[     346] = 32'hbcca629b;
    ram_cell[     347] = 32'ha0cf62fa;
    ram_cell[     348] = 32'h07898642;
    ram_cell[     349] = 32'hb5117049;
    ram_cell[     350] = 32'hf9574bf2;
    ram_cell[     351] = 32'h3c1439b1;
    ram_cell[     352] = 32'h06349740;
    ram_cell[     353] = 32'h40a1ccf0;
    ram_cell[     354] = 32'h4bfb1a91;
    ram_cell[     355] = 32'h5afb1695;
    ram_cell[     356] = 32'h458a0b4f;
    ram_cell[     357] = 32'h4dee6077;
    ram_cell[     358] = 32'hd631075f;
    ram_cell[     359] = 32'hac97b443;
    ram_cell[     360] = 32'hb6a103cf;
    ram_cell[     361] = 32'h9d8767e7;
    ram_cell[     362] = 32'h528ef0fc;
    ram_cell[     363] = 32'h0f5b4056;
    ram_cell[     364] = 32'hfece4390;
    ram_cell[     365] = 32'h7e080c09;
    ram_cell[     366] = 32'hafff8ec1;
    ram_cell[     367] = 32'h9494cbcc;
    ram_cell[     368] = 32'h78d3e4a4;
    ram_cell[     369] = 32'h9cee5323;
    ram_cell[     370] = 32'h09f6f2ef;
    ram_cell[     371] = 32'h21a7bc0b;
    ram_cell[     372] = 32'h24b1ab2a;
    ram_cell[     373] = 32'h61be469f;
    ram_cell[     374] = 32'he48be168;
    ram_cell[     375] = 32'h87ad82d2;
    ram_cell[     376] = 32'h3c2bb3bb;
    ram_cell[     377] = 32'he98a852a;
    ram_cell[     378] = 32'h5105fe3b;
    ram_cell[     379] = 32'h8d051e9a;
    ram_cell[     380] = 32'hf6b2a08c;
    ram_cell[     381] = 32'hab99141d;
    ram_cell[     382] = 32'h390a6efb;
    ram_cell[     383] = 32'hf99740a1;
    ram_cell[     384] = 32'h2a776839;
    ram_cell[     385] = 32'h5fa218e1;
    ram_cell[     386] = 32'h64b1e45c;
    ram_cell[     387] = 32'h2fb71e79;
    ram_cell[     388] = 32'hdc57aded;
    ram_cell[     389] = 32'h2c70a7ee;
    ram_cell[     390] = 32'h8a57c329;
    ram_cell[     391] = 32'hc1b0ed95;
    ram_cell[     392] = 32'hd01e139e;
    ram_cell[     393] = 32'ha5e364e3;
    ram_cell[     394] = 32'h9a36fbf9;
    ram_cell[     395] = 32'h06e531a6;
    ram_cell[     396] = 32'h5af7d672;
    ram_cell[     397] = 32'hb6cb2f0a;
    ram_cell[     398] = 32'h45acbc88;
    ram_cell[     399] = 32'hfe442bcf;
    ram_cell[     400] = 32'h2ef96dc7;
    ram_cell[     401] = 32'hbfa28f02;
    ram_cell[     402] = 32'hfd961721;
    ram_cell[     403] = 32'h08d129a0;
    ram_cell[     404] = 32'h1e67ba41;
    ram_cell[     405] = 32'he66610ca;
    ram_cell[     406] = 32'he89aa746;
    ram_cell[     407] = 32'h90df5ee1;
    ram_cell[     408] = 32'hd7d1c3a4;
    ram_cell[     409] = 32'h3cd73e6c;
    ram_cell[     410] = 32'h764b6d7a;
    ram_cell[     411] = 32'hc7b74b16;
    ram_cell[     412] = 32'hd508923b;
    ram_cell[     413] = 32'ha611fdfe;
    ram_cell[     414] = 32'hdc6d8525;
    ram_cell[     415] = 32'hf2037413;
    ram_cell[     416] = 32'h9872e039;
    ram_cell[     417] = 32'h8d911348;
    ram_cell[     418] = 32'h5284b129;
    ram_cell[     419] = 32'hdc1dbfe1;
    ram_cell[     420] = 32'h8c13abf9;
    ram_cell[     421] = 32'hc2328f81;
    ram_cell[     422] = 32'h1bfcf3af;
    ram_cell[     423] = 32'h2bc6570b;
    ram_cell[     424] = 32'h3a8aeed7;
    ram_cell[     425] = 32'h12dd3411;
    ram_cell[     426] = 32'h3ca20184;
    ram_cell[     427] = 32'h896c7ea8;
    ram_cell[     428] = 32'hf5f0aa8f;
    ram_cell[     429] = 32'h98aadef7;
    ram_cell[     430] = 32'hb46eef5e;
    ram_cell[     431] = 32'hbc534913;
    ram_cell[     432] = 32'hd4c9c27a;
    ram_cell[     433] = 32'h3eb07b90;
    ram_cell[     434] = 32'h4819b72f;
    ram_cell[     435] = 32'h99497fba;
    ram_cell[     436] = 32'h399ae219;
    ram_cell[     437] = 32'hd7c32cb2;
    ram_cell[     438] = 32'h73bf64b6;
    ram_cell[     439] = 32'h493d3f68;
    ram_cell[     440] = 32'hbd411c64;
    ram_cell[     441] = 32'hfc8617ad;
    ram_cell[     442] = 32'ha9a6565f;
    ram_cell[     443] = 32'hd31d01a2;
    ram_cell[     444] = 32'h29ff5198;
    ram_cell[     445] = 32'h76581bad;
    ram_cell[     446] = 32'h264f8439;
    ram_cell[     447] = 32'h55158d0a;
    ram_cell[     448] = 32'hd7300e92;
    ram_cell[     449] = 32'h559ce735;
    ram_cell[     450] = 32'hbe4c3549;
    ram_cell[     451] = 32'h755d8208;
    ram_cell[     452] = 32'hc267d8ec;
    ram_cell[     453] = 32'h94608b00;
    ram_cell[     454] = 32'h717ab834;
    ram_cell[     455] = 32'h0028a092;
    ram_cell[     456] = 32'h906c0589;
    ram_cell[     457] = 32'h60c60367;
    ram_cell[     458] = 32'h1a5d61e5;
    ram_cell[     459] = 32'h3ac5f3b2;
    ram_cell[     460] = 32'h26b2554a;
    ram_cell[     461] = 32'h7116729f;
    ram_cell[     462] = 32'h3d9cb3bb;
    ram_cell[     463] = 32'h62388407;
    ram_cell[     464] = 32'h778bf90d;
    ram_cell[     465] = 32'h76aa7f21;
    ram_cell[     466] = 32'hf334f5af;
    ram_cell[     467] = 32'h5259e3c3;
    ram_cell[     468] = 32'h00663a36;
    ram_cell[     469] = 32'h4dc2f016;
    ram_cell[     470] = 32'he5241f9e;
    ram_cell[     471] = 32'h1e5d35d7;
    ram_cell[     472] = 32'ha5570615;
    ram_cell[     473] = 32'h6ff151fd;
    ram_cell[     474] = 32'h93f12aac;
    ram_cell[     475] = 32'hbd4028f6;
    ram_cell[     476] = 32'h1401d435;
    ram_cell[     477] = 32'hff57ba5e;
    ram_cell[     478] = 32'hf23fdab6;
    ram_cell[     479] = 32'h8b26f874;
    ram_cell[     480] = 32'h270b86c0;
    ram_cell[     481] = 32'h430ff576;
    ram_cell[     482] = 32'h6f47c731;
    ram_cell[     483] = 32'h5d304ab7;
    ram_cell[     484] = 32'he9c49962;
    ram_cell[     485] = 32'h21f5d5f3;
    ram_cell[     486] = 32'ha06a8240;
    ram_cell[     487] = 32'h27e4a8a0;
    ram_cell[     488] = 32'h24edc466;
    ram_cell[     489] = 32'h98145bb8;
    ram_cell[     490] = 32'h67a0b987;
    ram_cell[     491] = 32'hae0a9aed;
    ram_cell[     492] = 32'hf5541d56;
    ram_cell[     493] = 32'heeb95062;
    ram_cell[     494] = 32'he91a27de;
    ram_cell[     495] = 32'hdbdd509e;
    ram_cell[     496] = 32'h75026bb5;
    ram_cell[     497] = 32'h767576b1;
    ram_cell[     498] = 32'ha0025710;
    ram_cell[     499] = 32'he8fa42a4;
    ram_cell[     500] = 32'hefef6253;
    ram_cell[     501] = 32'h166c92cb;
    ram_cell[     502] = 32'h8a5400c6;
    ram_cell[     503] = 32'h7dd477de;
    ram_cell[     504] = 32'hd284defd;
    ram_cell[     505] = 32'h2c77d66c;
    ram_cell[     506] = 32'h09c4f1f4;
    ram_cell[     507] = 32'h4d619033;
    ram_cell[     508] = 32'hf7c7077f;
    ram_cell[     509] = 32'h2709c48c;
    ram_cell[     510] = 32'h0d0935f0;
    ram_cell[     511] = 32'h3e9d1638;
    // src matrix B
    ram_cell[     512] = 32'h095ee730;
    ram_cell[     513] = 32'h7d0c4ae7;
    ram_cell[     514] = 32'h924cb44e;
    ram_cell[     515] = 32'ha24cf1fd;
    ram_cell[     516] = 32'h1642c48c;
    ram_cell[     517] = 32'hfb6b6ab8;
    ram_cell[     518] = 32'he257055d;
    ram_cell[     519] = 32'hcc94e53d;
    ram_cell[     520] = 32'hfdf02e97;
    ram_cell[     521] = 32'had6d96bb;
    ram_cell[     522] = 32'h81ea7368;
    ram_cell[     523] = 32'he3c23abd;
    ram_cell[     524] = 32'h0bece69e;
    ram_cell[     525] = 32'hce3d7c38;
    ram_cell[     526] = 32'h0d01d395;
    ram_cell[     527] = 32'hac2d1d10;
    ram_cell[     528] = 32'h2a577515;
    ram_cell[     529] = 32'h132ce1cb;
    ram_cell[     530] = 32'h0c1d7381;
    ram_cell[     531] = 32'h62b94714;
    ram_cell[     532] = 32'h349af6e9;
    ram_cell[     533] = 32'h5e9dced7;
    ram_cell[     534] = 32'ha67e3e03;
    ram_cell[     535] = 32'he0b979fb;
    ram_cell[     536] = 32'h09905ba1;
    ram_cell[     537] = 32'had17e9a1;
    ram_cell[     538] = 32'hab37e2af;
    ram_cell[     539] = 32'ha758cbfd;
    ram_cell[     540] = 32'h086eaacf;
    ram_cell[     541] = 32'hf8232071;
    ram_cell[     542] = 32'hc7058fb7;
    ram_cell[     543] = 32'h31af9dfe;
    ram_cell[     544] = 32'h807bf118;
    ram_cell[     545] = 32'h6cb52c95;
    ram_cell[     546] = 32'hc039649e;
    ram_cell[     547] = 32'hc46f87e6;
    ram_cell[     548] = 32'hac3b79dc;
    ram_cell[     549] = 32'hd7399821;
    ram_cell[     550] = 32'h1eadca2a;
    ram_cell[     551] = 32'hbb5b0e25;
    ram_cell[     552] = 32'h15c53b7c;
    ram_cell[     553] = 32'hada909ca;
    ram_cell[     554] = 32'h65488808;
    ram_cell[     555] = 32'h8c94c97f;
    ram_cell[     556] = 32'ha26be745;
    ram_cell[     557] = 32'h9d969301;
    ram_cell[     558] = 32'h601a1890;
    ram_cell[     559] = 32'h2e1367f0;
    ram_cell[     560] = 32'h20909187;
    ram_cell[     561] = 32'h44a26bea;
    ram_cell[     562] = 32'h8e3f6407;
    ram_cell[     563] = 32'h1b57c65f;
    ram_cell[     564] = 32'h664c9b0f;
    ram_cell[     565] = 32'haf7ec129;
    ram_cell[     566] = 32'h0509d1aa;
    ram_cell[     567] = 32'h94565808;
    ram_cell[     568] = 32'h6cb39d50;
    ram_cell[     569] = 32'h5088868c;
    ram_cell[     570] = 32'h0ed2ae92;
    ram_cell[     571] = 32'ha52b0ab9;
    ram_cell[     572] = 32'h6cd4cb31;
    ram_cell[     573] = 32'hcbf2c493;
    ram_cell[     574] = 32'h3e2e6540;
    ram_cell[     575] = 32'h80274508;
    ram_cell[     576] = 32'h3607e4e4;
    ram_cell[     577] = 32'haa43bc2b;
    ram_cell[     578] = 32'hff0131d2;
    ram_cell[     579] = 32'hdea70ccf;
    ram_cell[     580] = 32'h8ca9dfd2;
    ram_cell[     581] = 32'hd783b930;
    ram_cell[     582] = 32'h3035f19b;
    ram_cell[     583] = 32'he3da1d14;
    ram_cell[     584] = 32'h4842a9ab;
    ram_cell[     585] = 32'h791cbe0b;
    ram_cell[     586] = 32'h201bf167;
    ram_cell[     587] = 32'h1ea264b5;
    ram_cell[     588] = 32'he444ec23;
    ram_cell[     589] = 32'h4dd1adb2;
    ram_cell[     590] = 32'h210ff608;
    ram_cell[     591] = 32'hc24a163a;
    ram_cell[     592] = 32'he31ff360;
    ram_cell[     593] = 32'hdb851c07;
    ram_cell[     594] = 32'hce099504;
    ram_cell[     595] = 32'hc546723d;
    ram_cell[     596] = 32'h88040fc6;
    ram_cell[     597] = 32'h468f530d;
    ram_cell[     598] = 32'hd727d312;
    ram_cell[     599] = 32'h44c0373b;
    ram_cell[     600] = 32'hdb17fae3;
    ram_cell[     601] = 32'h758730a2;
    ram_cell[     602] = 32'h34450aad;
    ram_cell[     603] = 32'h928d398e;
    ram_cell[     604] = 32'h0454e33f;
    ram_cell[     605] = 32'haf7e41ed;
    ram_cell[     606] = 32'h2d95a2e3;
    ram_cell[     607] = 32'h15258cee;
    ram_cell[     608] = 32'h42a8c53b;
    ram_cell[     609] = 32'h0d09c6c6;
    ram_cell[     610] = 32'hdf016553;
    ram_cell[     611] = 32'he7d47877;
    ram_cell[     612] = 32'ha60429b3;
    ram_cell[     613] = 32'hc40e1602;
    ram_cell[     614] = 32'hf0ac1614;
    ram_cell[     615] = 32'h4ff059a9;
    ram_cell[     616] = 32'h8f377278;
    ram_cell[     617] = 32'hcee07e8d;
    ram_cell[     618] = 32'hecde8b94;
    ram_cell[     619] = 32'h0be9912e;
    ram_cell[     620] = 32'hb258d714;
    ram_cell[     621] = 32'h52b7acb8;
    ram_cell[     622] = 32'h1ad6e40b;
    ram_cell[     623] = 32'hc690c767;
    ram_cell[     624] = 32'h0a32d1a9;
    ram_cell[     625] = 32'h5a60dcc9;
    ram_cell[     626] = 32'h6736c9d2;
    ram_cell[     627] = 32'ha2914a4e;
    ram_cell[     628] = 32'hf1c49ed8;
    ram_cell[     629] = 32'hef230d80;
    ram_cell[     630] = 32'ha9f79859;
    ram_cell[     631] = 32'h56a10202;
    ram_cell[     632] = 32'h0c6d5ddc;
    ram_cell[     633] = 32'h47243e30;
    ram_cell[     634] = 32'haa753c0a;
    ram_cell[     635] = 32'hbebb8acb;
    ram_cell[     636] = 32'h0918652b;
    ram_cell[     637] = 32'h166c7796;
    ram_cell[     638] = 32'h132061e9;
    ram_cell[     639] = 32'hc1e738bb;
    ram_cell[     640] = 32'h89b16bf3;
    ram_cell[     641] = 32'h07145724;
    ram_cell[     642] = 32'hb3daa000;
    ram_cell[     643] = 32'h099d8dc3;
    ram_cell[     644] = 32'h73e15226;
    ram_cell[     645] = 32'h73d3157c;
    ram_cell[     646] = 32'h4b149c4d;
    ram_cell[     647] = 32'hd917aa17;
    ram_cell[     648] = 32'h54b79218;
    ram_cell[     649] = 32'h8c468b69;
    ram_cell[     650] = 32'hb9ab9a3f;
    ram_cell[     651] = 32'hcb25243b;
    ram_cell[     652] = 32'h94fed73b;
    ram_cell[     653] = 32'hde39278a;
    ram_cell[     654] = 32'h9d57325f;
    ram_cell[     655] = 32'h648b3d71;
    ram_cell[     656] = 32'h19d29f8a;
    ram_cell[     657] = 32'h97d239c0;
    ram_cell[     658] = 32'h4c285656;
    ram_cell[     659] = 32'h641f13a8;
    ram_cell[     660] = 32'h97ad25ba;
    ram_cell[     661] = 32'h1666090b;
    ram_cell[     662] = 32'h104f0455;
    ram_cell[     663] = 32'hca6dfc59;
    ram_cell[     664] = 32'h74b432a4;
    ram_cell[     665] = 32'h28987fdf;
    ram_cell[     666] = 32'hc76905d8;
    ram_cell[     667] = 32'hd4c48cc7;
    ram_cell[     668] = 32'h8d9da730;
    ram_cell[     669] = 32'hb94742d0;
    ram_cell[     670] = 32'h81d11fc9;
    ram_cell[     671] = 32'h51be735c;
    ram_cell[     672] = 32'hf8e94d0c;
    ram_cell[     673] = 32'hf2a4a634;
    ram_cell[     674] = 32'hc3534120;
    ram_cell[     675] = 32'h6550267c;
    ram_cell[     676] = 32'h9fc51a8f;
    ram_cell[     677] = 32'ha1947e9a;
    ram_cell[     678] = 32'hfa7dbf7d;
    ram_cell[     679] = 32'h0d8c000b;
    ram_cell[     680] = 32'h0e68c75d;
    ram_cell[     681] = 32'h1602fbec;
    ram_cell[     682] = 32'h8c638b2c;
    ram_cell[     683] = 32'he9350f32;
    ram_cell[     684] = 32'h5efe3aa2;
    ram_cell[     685] = 32'h58f5b0f2;
    ram_cell[     686] = 32'h8aa6147a;
    ram_cell[     687] = 32'hfaafa1eb;
    ram_cell[     688] = 32'h28ae93e5;
    ram_cell[     689] = 32'h3c9e7f07;
    ram_cell[     690] = 32'h57ef9dc4;
    ram_cell[     691] = 32'hb5350b99;
    ram_cell[     692] = 32'h9c4f30d3;
    ram_cell[     693] = 32'hb1a61c56;
    ram_cell[     694] = 32'hb21466a6;
    ram_cell[     695] = 32'hb26d4436;
    ram_cell[     696] = 32'hd0bdf8a2;
    ram_cell[     697] = 32'h5b803890;
    ram_cell[     698] = 32'h73deb2d1;
    ram_cell[     699] = 32'hcc4afb02;
    ram_cell[     700] = 32'h2aec4b2e;
    ram_cell[     701] = 32'h2bf0ff1f;
    ram_cell[     702] = 32'h758bee32;
    ram_cell[     703] = 32'hed33e26b;
    ram_cell[     704] = 32'h0bc3b480;
    ram_cell[     705] = 32'hf87189df;
    ram_cell[     706] = 32'h084212c2;
    ram_cell[     707] = 32'h37a7a31e;
    ram_cell[     708] = 32'h7e4f7504;
    ram_cell[     709] = 32'h2f83ab05;
    ram_cell[     710] = 32'h1842834a;
    ram_cell[     711] = 32'h944b5311;
    ram_cell[     712] = 32'ha03e23dc;
    ram_cell[     713] = 32'h5640683a;
    ram_cell[     714] = 32'h1dd2d1cb;
    ram_cell[     715] = 32'hc3b93fb5;
    ram_cell[     716] = 32'hfe5c3459;
    ram_cell[     717] = 32'h3e7c9fed;
    ram_cell[     718] = 32'h6d4a51bd;
    ram_cell[     719] = 32'he27251ad;
    ram_cell[     720] = 32'hfc31281d;
    ram_cell[     721] = 32'h28198646;
    ram_cell[     722] = 32'h122271a3;
    ram_cell[     723] = 32'h75bc2fe5;
    ram_cell[     724] = 32'he427d1ef;
    ram_cell[     725] = 32'hf7d87662;
    ram_cell[     726] = 32'h6007e29f;
    ram_cell[     727] = 32'h036e346f;
    ram_cell[     728] = 32'hb06708da;
    ram_cell[     729] = 32'h501dfc19;
    ram_cell[     730] = 32'hb12a32ca;
    ram_cell[     731] = 32'hdbcb725a;
    ram_cell[     732] = 32'h87d84726;
    ram_cell[     733] = 32'hc156b490;
    ram_cell[     734] = 32'h7b4274de;
    ram_cell[     735] = 32'h4038797f;
    ram_cell[     736] = 32'h7369e7a6;
    ram_cell[     737] = 32'ha7a99b5e;
    ram_cell[     738] = 32'hac234c9f;
    ram_cell[     739] = 32'h0034f924;
    ram_cell[     740] = 32'hb24cf500;
    ram_cell[     741] = 32'h70ac8808;
    ram_cell[     742] = 32'h36a4f67f;
    ram_cell[     743] = 32'h94b975f7;
    ram_cell[     744] = 32'h0cefef37;
    ram_cell[     745] = 32'h605c006a;
    ram_cell[     746] = 32'he478122e;
    ram_cell[     747] = 32'h8533eeda;
    ram_cell[     748] = 32'h29b4b97a;
    ram_cell[     749] = 32'h3a97f5fa;
    ram_cell[     750] = 32'h381ec1ba;
    ram_cell[     751] = 32'h0373b4da;
    ram_cell[     752] = 32'h208d0231;
    ram_cell[     753] = 32'h3fcd7400;
    ram_cell[     754] = 32'h7789008d;
    ram_cell[     755] = 32'h4cff6e46;
    ram_cell[     756] = 32'hfb763378;
    ram_cell[     757] = 32'hd09c9fb1;
    ram_cell[     758] = 32'h91ec5b28;
    ram_cell[     759] = 32'h65584653;
    ram_cell[     760] = 32'h2485be75;
    ram_cell[     761] = 32'h88a4dc1e;
    ram_cell[     762] = 32'hdb3482ab;
    ram_cell[     763] = 32'h1ef8f02e;
    ram_cell[     764] = 32'ha303cdd6;
    ram_cell[     765] = 32'h3c46b28a;
    ram_cell[     766] = 32'h081f8561;
    ram_cell[     767] = 32'h47c2e352;
end

endmodule

